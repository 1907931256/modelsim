timescale 1 ns/1 ps
module PCI_LC_I (
  OE_DEVSEL, BASE_HIT0, BASE_HIT1, BASE_HIT2, BASE_HIT3, BASE_HIT4, BASE_HIT5, BASE_HIT6, BASE_HIT7, S_DATA_VLD, OE_REQ, OE_CBE, OE_ADO_LT64, OE_IRDY
, REQUEST64, SLOT64, IRDY_I, IRDY_O, AD10, AD11, AD12, AD13, AD14, AD15, AD16, AD0, AD17, AD20, AD1, AD18, AD21, AD2, AD19, AD22, AD3, AD23, AD4, AD24
, AD5, AD25, AD6, AD26, AD7, AD27, AD30, AD8, AD28, AD31, AD9, AD29, AD32, AD33, CSR10, AD34, PAR64_I, CSR11, CLKX, AD35, CSR12, AD36, M_ADDR_N, CSR13
, AD37, CSR14, AD40, AD38, CSR15, AD41, AD39, CSR16, AD42, AD_O10, PAR64_O, CSR20, CSR17, AD43, AD_O11, CSR21, CSR18, AD44, AD_O12, CSR22, CSR19, AD45
, AD_O13, CSR23, ACK64_I, AD46, AD_O14, CSR24, AD47, AD50, AD_O15, CSR25, AD48, AD51, AD_O16, CSR26, AD49, AD52, AD_O17, CSR30, CSR27, AD_O20, AD53, 
AD_O18, CSR31, CSR28, AD_O21, AD54, AD_O19, CSR32, CSR29, AD_O22, ACK64_O, AD55, AD_O23, CSR33, AD56, AD_O24, CSR34, AD57, AD60, AD_O25, CSR35, AD58, 
AD61, AD_O26, CSR36, AD59, AD62, AD_O27, CSR37, AD_O30, AD63, AD_O28, CSR38, AD_O31, AD_O29, CSR39, AD_O32, AD_O33, AD_O34, AD_O35, AD_O36, AD_O40, 
AD_O37, AD_O41, AD_O38, AD_O42, AD_O39, AD_O43, AD_O44, AD_O45, AD_O46, AD_O50, AD_O47, AD_O51, AD_O48, AD_O52, SERRQ_N, AD_O49, AD_O53, AD_O54, 
AD_O55, AD_O56, PAR_I, AD_O60, AD_O57, ADIO0, AD_O61, AD_O58, ADIO1, AD_O62, AD_O59, ADIO2, AD_O63, ADIO3, STOP_I, ADIO4, PAR_O, ADIO5, ADIO6, ADIO7, 
S_CYCLE64, ADIO8, ADIO9, STOP_O, S_SRC_EN, PERRQ_N, M_CBE0, M_CBE1, M_CBE2, M_CBE3, M_CBE4, M_CBE5, M_CBE6, M_CBE7, M_WRDN, PERR_I, CBE_IN0, CBE_IN1, 
CBE_IN2, PERR_O, CBE_IN3, INTR_N, CBE_IN4, CBE_IN5, CBE_IN6, CBE_IN7, CFG_SELF, IDLE, S_READY, DR_BUS, REQ64Q_N, PCI_CMD0, PCI_CMD1, PCI_CMD2, 
PCI_CMD3, PCI_CMD4, PCI_CMD5, PCI_CMD6, PCI_CMD7, PCI_CMD8, PCI_CMD9, S_TERM, IDSEL_IN, M_READY, COMPLETE, FRAME_I, S_CBE0, S_CBE1, S_CBE2, S_CBE3, 
ADDR_VLD, S_CBE4, FRAME_O, S_CBE5, S_CBE6, S_CBE7, S_WRDN, CLK, M_DATA_VLD, REQ64_I, OE_PERR, REQ64_O, RST, ACK64Q_N, GNT_IN, M_FAIL64, C_READY, 
PCI_CMD10, PCI_CMD11, PCI_CMD12, PCI_CMD13, PCI_CMD14, PCI_CMD15, TRDY_I, TRDY_O, OE_ACK64, DEVSELQ_N, CSR0, AD_O0, CSR1, AD_O1, CSR2, AD_O2, CSR3, 
AD_O3, CSR4, AD_O4, CSR5, AD_O5, CSR6, AD_O6, CSR7, AD_O7, CSR8, AD_O8, CSR9, AD_O9, ADDR10, ADDR11, ADDR12, ADDR13, ADDR14, ADDR15, ADDR16, ADDR20, 
ADDR17, ADDR21, ADDR18, ADDR22, ADDR19, ADDR23, ADDR24, ADDR25, ADDR26, ADDR30, ADDR27, ADDR31, ADDR28, ADDR29, DEVSEL_I, RST_N, DEVSEL_O, ADIO10, 
ADIO11, ADIO12, ADIO13, ADIO14, ADIO15, ADIO16, ADIO20, ADIO17, ADIO21, ADIO18, ADIO22, ADIO19, ADIO23, ADIO24, ADIO25, ADIO26, ADIO30, ADIO27, ADIO31
, ADIO28, CFG0, ADIO32, ADIO29, CFG1, ADIO33, CFG2, ADIO34, CFG3, ADIO35, CFG4, ADIO36, CFG5, ADIO37, CFG6, ADIO40, ADIO38, CFG7, ADIO41, ADIO39, CFG8
, ADIO42, CFG10, CFG9, ADIO43, CFG11, ADIO44, CFG12, ADIO45, CFG13, ADIO46, CFG14, ADIO47, ADIO50, CFG15, ADIO48, ADIO51, CFG16, ADIO49, ADIO52, CFG17
, C_TERM, CFG20, ADIO53, CFG18, OE_ADO_B, CFG21, ADIO54, CFG19, CFG22, ADIO55, ADIO56, CFG23, ADIO57, M_SRC_EN, CFG24, ADIO60, ADIO58, CFG25, ADIO61, 
ADIO59, CFG26, ADIO62, ADIO63, CFG30, CFG27, CFG28, CFG31, CFG29, CFG32, CFG33, CFG34, CFG35, CFG36, CFG37, CFG40, CFG38, CFG41, CFG39, CFG42, CFG43, 
CFG44, CFG45, OE_ADO_T, CFG46, CFG47, CFG50, CFG48, CFG51, CFG49, CFG52, CFG53, CFG54, SUB_DATA10, REQ_OUT, CFG55, SUB_DATA11, CFG56, SUB_DATA12, 
CFG57, SUB_DATA13, CFG60, CFG58, SUB_DATA14, CFG61, CFG59, SUB_DATA15, CFG62, CFG63, SUB_DATA16, CFG64, SUB_DATA20, SUB_DATA17, CFG65, SUB_DATA21, 
SUB_DATA18, OE_STOP, CFG66, SUB_DATA22, SUB_DATA19, CFG67, SUB_DATA23, CFG70, CFG68, SUB_DATA24, CFG71, CFG69, SUB_DATA25, CFG72, CFG73, SUB_DATA26, 
CFG74, SUB_DATA30, SUB_DATA27, CFG75, SUB_DATA31, SUB_DATA28, CFG76, SUB_DATA29, CFG77, CFG80, CFG78, CFG81, CFG79, TIME_OUT, CFG82, CFG83, CFG84, 
CFG85, CFG86, TRDYQ_N, CFG100, CFG90, CFG87, CFG101, CFG91, CFG88, CFG102, CFG92, CFG89, CFG103, CFG93, CFG104, CFG94, CFG105, CFG95, CFG106, CFG96, 
CFG107, CFG97, CFG110, CFG108, CFG98, CFG111, CFG109, CFG99, CFG112, CFG113, CFG114, CFG115, CFG116, CFG117, CFG120, CFG118, CFG121, CFG119, CFG122, 
CFG123, CFG124, CFG125, CFG126, CFG127, CFG130, CFG128, CFG131, CFG129, CFG132, CFG133, CFG134, OE_FRAME, CFG135, CFG136, I_IDLE, CFG137, CFG140, 
CFG138, CFG141, CFG139, CFG142, CFG143, CFG144, CFG145, CFG146, CFG147, CFG150, CFG148, CFG151, CFG149, CFG152, CFG153, CFG154, STOPQ_N, CFG155, 
CFG156, OE_SERR, CFG157, OE_ADO_B64, CFG160, CFG158, CFG161, CFG159, CFG162, CFG163, CFG164, CFG165, CFG166, CFG170, CFG200, CFG167, CFG171, CFG201, 
CFG168, CFG172, CFG202, CFG169, CFG203, CFG173, CBE_I0, CFG204, CFG174, CBE_I1, CFG175, CFG205, CBE_I2, CFG206, CFG176, CBE_I3, CFG180, CFG207, CFG210
, CFG177, CBE_I4, CFG181, CFG208, CFG211, CFG178, CBE_I5, CFG212, CFG182, CFG209, CFG179, CBE_I6, CFG213, CFG183, CBE_I7, CFG214, CFG184, CFG185, 
CFG215, CFG186, CFG216, CFG190, CFG220, CFG217, CFG187, CFG191, CFG221, CFG218, CFG188, CFG192, CFG222, CFG219, CFG189, CFG193, CFG223, CFG194, CFG224
, CFG195, CFG225, CFG196, CFG226, CFG197, CFG230, CFG227, CFG198, CFG231, CFG228, CFG199, CFG232, CFG229, CFG233, B_BUSY, CFG234, CFG235, CFG236, 
CFG237, CFG240, CFG238, CFG_VLD, CFG241, CFG239, CFG242, CFG243, M_DATA, CFG244, CFG245, CFG246, CFG247, CFG250, CFG248, CFG251, CFG249, CFG252, 
CFG253, IRDYQ_N, CFG254, CFG255, SERR_I, CBE_O0, OE_PAR, CBE_O1, CBE_O2, REQUEST, CBE_O3, CBE_O4, CBE_O5, CBE_O6, CBE_O7, OE_ADO_LB64, OE_REQ64, 
KEEPOUT, OE_INTA, REQUESTHOLD, S_ABORT, ADDR0, OE_PAR64, ADDR1, ADDR2, ADDR3, ADDR4, ADDR5, ADDR6, BACKOFF, ADDR7, ADDR8, OE_ADO_T64, ADDR9, CFG_HIT, 
OE_TRDY, SUB_DATA0, SUB_DATA1, SUB_DATA2, SUB_DATA3, SUB_DATA4, SUB_DATA5, SUB_DATA6, OE_CBE64, SUB_DATA7, SUB_DATA8, SUB_DATA9, FRAMEQ_N, OE_ADO_LB, 
S_DATA, OE_ADO_LT
);
// synthesis attribute syn_edif_bit_format = "%u<%i>"
// synthesis attribute syn_edif_scalar_format = "%u"
// synthesis attribute syn_noclockbuf = 1
// synthesis attribute syn_hier = "hard"
// synthesis attribute syn_black_box
  output OE_DEVSEL;
  output BASE_HIT0;
  output BASE_HIT1;
  output BASE_HIT2;
  output BASE_HIT3;
  output BASE_HIT4;
  output BASE_HIT5;
  output BASE_HIT6;
  output BASE_HIT7;
  output S_DATA_VLD;
  output OE_REQ;
  output OE_CBE;
  output OE_ADO_LT64;
  output OE_IRDY;
  input REQUEST64;
  input SLOT64;
  input IRDY_I;
  output IRDY_O;
  input AD10;
  input AD11;
  input AD12;
  input AD13;
  input AD14;
  input AD15;
  input AD16;
  input AD0;
  input AD17;
  input AD20;
  input AD1;
  input AD18;
  input AD21;
  input AD2;
  input AD19;
  input AD22;
  input AD3;
  input AD23;
  input AD4;
  input AD24;
  input AD5;
  input AD25;
  input AD6;
  input AD26;
  input AD7;
  input AD27;
  input AD30;
  input AD8;
  input AD28;
  input AD31;
  input AD9;
  input AD29;
  input AD32;
  input AD33;
  output CSR10;
  input AD34;
  input PAR64_I;
  output CSR11;
  input CLKX;
  input AD35;
  output CSR12;
  input AD36;
  output M_ADDR_N;
  output CSR13;
  input AD37;
  output CSR14;
  input AD40;
  input AD38;
  output CSR15;
  input AD41;
  input AD39;
  output CSR16;
  input AD42;
  output AD_O10;
  output PAR64_O;
  output CSR20;
  output CSR17;
  input AD43;
  output AD_O11;
  output CSR21;
  output CSR18;
  input AD44;
  output AD_O12;
  output CSR22;
  output CSR19;
  input AD45;
  output AD_O13;
  output CSR23;
  input ACK64_I;
  input AD46;
  output AD_O14;
  output CSR24;
  input AD47;
  input AD50;
  output AD_O15;
  output CSR25;
  input AD48;
  input AD51;
  output AD_O16;
  output CSR26;
  input AD49;
  input AD52;
  output AD_O17;
  output CSR30;
  output CSR27;
  output AD_O20;
  input AD53;
  output AD_O18;
  output CSR31;
  output CSR28;
  output AD_O21;
  input AD54;
  output AD_O19;
  output CSR32;
  output CSR29;
  output AD_O22;
  output ACK64_O;
  input AD55;
  output AD_O23;
  output CSR33;
  input AD56;
  output AD_O24;
  output CSR34;
  input AD57;
  input AD60;
  output AD_O25;
  output CSR35;
  input AD58;
  input AD61;
  output AD_O26;
  output CSR36;
  input AD59;
  input AD62;
  output AD_O27;
  output CSR37;
  output AD_O30;
  input AD63;
  output AD_O28;
  output CSR38;
  output AD_O31;
  output AD_O29;
  output CSR39;
  output AD_O32;
  output AD_O33;
  output AD_O34;
  output AD_O35;
  output AD_O36;
  output AD_O40;
  output AD_O37;
  output AD_O41;
  output AD_O38;
  output AD_O42;
  output AD_O39;
  output AD_O43;
  output AD_O44;
  output AD_O45;
  output AD_O46;
  output AD_O50;
  output AD_O47;
  output AD_O51;
  output AD_O48;
  output AD_O52;
  output SERRQ_N;
  output AD_O49;
  output AD_O53;
  output AD_O54;
  output AD_O55;
  output AD_O56;
  input PAR_I;
  output AD_O60;
  output AD_O57;
  inout ADIO0;
  output AD_O61;
  output AD_O58;
  inout ADIO1;
  output AD_O62;
  output AD_O59;
  inout ADIO2;
  output AD_O63;
  inout ADIO3;
  input STOP_I;
  inout ADIO4;
  output PAR_O;
  inout ADIO5;
  inout ADIO6;
  inout ADIO7;
  output S_CYCLE64;
  inout ADIO8;
  inout ADIO9;
  output STOP_O;
  output S_SRC_EN;
  output PERRQ_N;
  input M_CBE0;
  input M_CBE1;
  input M_CBE2;
  input M_CBE3;
  input M_CBE4;
  input M_CBE5;
  input M_CBE6;
  input M_CBE7;
  input M_WRDN;
  input PERR_I;
  input CBE_IN0;
  input CBE_IN1;
  input CBE_IN2;
  output PERR_O;
  input CBE_IN3;
  input INTR_N;
  input CBE_IN4;
  input CBE_IN5;
  input CBE_IN6;
  input CBE_IN7;
  input CFG_SELF;
  output IDLE;
  input S_READY;
  output DR_BUS;
  output REQ64Q_N;
  output PCI_CMD0;
  output PCI_CMD1;
  output PCI_CMD2;
  output PCI_CMD3;
  output PCI_CMD4;
  output PCI_CMD5;
  output PCI_CMD6;
  output PCI_CMD7;
  output PCI_CMD8;
  output PCI_CMD9;
  input S_TERM;
  input IDSEL_IN;
  input M_READY;
  input COMPLETE;
  input FRAME_I;
  output S_CBE0;
  output S_CBE1;
  output S_CBE2;
  output S_CBE3;
  output ADDR_VLD;
  output S_CBE4;
  output FRAME_O;
  output S_CBE5;
  output S_CBE6;
  output S_CBE7;
  output S_WRDN;
  input CLK;
  output M_DATA_VLD;
  input REQ64_I;
  output OE_PERR;
  output REQ64_O;
  output RST;
  output ACK64Q_N;
  input GNT_IN;
  output M_FAIL64;
  input C_READY;
  output PCI_CMD10;
  output PCI_CMD11;
  output PCI_CMD12;
  output PCI_CMD13;
  output PCI_CMD14;
  output PCI_CMD15;
  input TRDY_I;
  output TRDY_O;
  output OE_ACK64;
  output DEVSELQ_N;
  output CSR0;
  output AD_O0;
  output CSR1;
  output AD_O1;
  output CSR2;
  output AD_O2;
  output CSR3;
  output AD_O3;
  output CSR4;
  output AD_O4;
  output CSR5;
  output AD_O5;
  output CSR6;
  output AD_O6;
  output CSR7;
  output AD_O7;
  output CSR8;
  output AD_O8;
  output CSR9;
  output AD_O9;
  output ADDR10;
  output ADDR11;
  output ADDR12;
  output ADDR13;
  output ADDR14;
  output ADDR15;
  output ADDR16;
  output ADDR20;
  output ADDR17;
  output ADDR21;
  output ADDR18;
  output ADDR22;
  output ADDR19;
  output ADDR23;
  output ADDR24;
  output ADDR25;
  output ADDR26;
  output ADDR30;
  output ADDR27;
  output ADDR31;
  output ADDR28;
  output ADDR29;
  input DEVSEL_I;
  input RST_N;
  output DEVSEL_O;
  inout ADIO10;
  inout ADIO11;
  inout ADIO12;
  inout ADIO13;
  inout ADIO14;
  inout ADIO15;
  inout ADIO16;
  inout ADIO20;
  inout ADIO17;
  inout ADIO21;
  inout ADIO18;
  inout ADIO22;
  inout ADIO19;
  inout ADIO23;
  inout ADIO24;
  inout ADIO25;
  inout ADIO26;
  inout ADIO30;
  inout ADIO27;
  inout ADIO31;
  inout ADIO28;
  input CFG0;
  inout ADIO32;
  inout ADIO29;
  input CFG1;
  inout ADIO33;
  input CFG2;
  inout ADIO34;
  input CFG3;
  inout ADIO35;
  input CFG4;
  inout ADIO36;
  input CFG5;
  inout ADIO37;
  input CFG6;
  inout ADIO40;
  inout ADIO38;
  input CFG7;
  inout ADIO41;
  inout ADIO39;
  input CFG8;
  inout ADIO42;
  input CFG10;
  input CFG9;
  inout ADIO43;
  input CFG11;
  inout ADIO44;
  input CFG12;
  inout ADIO45;
  input CFG13;
  inout ADIO46;
  input CFG14;
  inout ADIO47;
  inout ADIO50;
  input CFG15;
  inout ADIO48;
  inout ADIO51;
  input CFG16;
  inout ADIO49;
  inout ADIO52;
  input CFG17;
  input C_TERM;
  input CFG20;
  inout ADIO53;
  input CFG18;
  output OE_ADO_B;
  input CFG21;
  inout ADIO54;
  input CFG19;
  input CFG22;
  inout ADIO55;
  inout ADIO56;
  input CFG23;
  inout ADIO57;
  output M_SRC_EN;
  input CFG24;
  inout ADIO60;
  inout ADIO58;
  input CFG25;
  inout ADIO61;
  inout ADIO59;
  input CFG26;
  inout ADIO62;
  inout ADIO63;
  input CFG30;
  input CFG27;
  input CFG28;
  input CFG31;
  input CFG29;
  input CFG32;
  input CFG33;
  input CFG34;
  input CFG35;
  input CFG36;
  input CFG37;
  input CFG40;
  input CFG38;
  input CFG41;
  input CFG39;
  input CFG42;
  input CFG43;
  input CFG44;
  input CFG45;
  output OE_ADO_T;
  input CFG46;
  input CFG47;
  input CFG50;
  input CFG48;
  input CFG51;
  input CFG49;
  input CFG52;
  input CFG53;
  input CFG54;
  input SUB_DATA10;
  output REQ_OUT;
  input CFG55;
  input SUB_DATA11;
  input CFG56;
  input SUB_DATA12;
  input CFG57;
  input SUB_DATA13;
  input CFG60;
  input CFG58;
  input SUB_DATA14;
  input CFG61;
  input CFG59;
  input SUB_DATA15;
  input CFG62;
  input CFG63;
  input SUB_DATA16;
  input CFG64;
  input SUB_DATA20;
  input SUB_DATA17;
  input CFG65;
  input SUB_DATA21;
  input SUB_DATA18;
  output OE_STOP;
  input CFG66;
  input SUB_DATA22;
  input SUB_DATA19;
  input CFG67;
  input SUB_DATA23;
  input CFG70;
  input CFG68;
  input SUB_DATA24;
  input CFG71;
  input CFG69;
  input SUB_DATA25;
  input CFG72;
  input CFG73;
  input SUB_DATA26;
  input CFG74;
  input SUB_DATA30;
  input SUB_DATA27;
  input CFG75;
  input SUB_DATA31;
  input SUB_DATA28;
  input CFG76;
  input SUB_DATA29;
  input CFG77;
  input CFG80;
  input CFG78;
  input CFG81;
  input CFG79;
  output TIME_OUT;
  input CFG82;
  input CFG83;
  input CFG84;
  input CFG85;
  input CFG86;
  output TRDYQ_N;
  input CFG100;
  input CFG90;
  input CFG87;
  input CFG101;
  input CFG91;
  input CFG88;
  input CFG102;
  input CFG92;
  input CFG89;
  input CFG103;
  input CFG93;
  input CFG104;
  input CFG94;
  input CFG105;
  input CFG95;
  input CFG106;
  input CFG96;
  input CFG107;
  input CFG97;
  input CFG110;
  input CFG108;
  input CFG98;
  input CFG111;
  input CFG109;
  input CFG99;
  input CFG112;
  input CFG113;
  input CFG114;
  input CFG115;
  input CFG116;
  input CFG117;
  input CFG120;
  input CFG118;
  input CFG121;
  input CFG119;
  input CFG122;
  input CFG123;
  input CFG124;
  input CFG125;
  input CFG126;
  input CFG127;
  input CFG130;
  input CFG128;
  input CFG131;
  input CFG129;
  input CFG132;
  input CFG133;
  input CFG134;
  output OE_FRAME;
  input CFG135;
  input CFG136;
  output I_IDLE;
  input CFG137;
  input CFG140;
  input CFG138;
  input CFG141;
  input CFG139;
  input CFG142;
  input CFG143;
  input CFG144;
  input CFG145;
  input CFG146;
  input CFG147;
  input CFG150;
  input CFG148;
  input CFG151;
  input CFG149;
  input CFG152;
  input CFG153;
  input CFG154;
  output STOPQ_N;
  input CFG155;
  input CFG156;
  output OE_SERR;
  input CFG157;
  output OE_ADO_B64;
  input CFG160;
  input CFG158;
  input CFG161;
  input CFG159;
  input CFG162;
  input CFG163;
  input CFG164;
  input CFG165;
  input CFG166;
  input CFG170;
  input CFG200;
  input CFG167;
  input CFG171;
  input CFG201;
  input CFG168;
  input CFG172;
  input CFG202;
  input CFG169;
  input CFG203;
  input CFG173;
  input CBE_I0;
  input CFG204;
  input CFG174;
  input CBE_I1;
  input CFG175;
  input CFG205;
  input CBE_I2;
  input CFG206;
  input CFG176;
  input CBE_I3;
  input CFG180;
  input CFG207;
  input CFG210;
  input CFG177;
  input CBE_I4;
  input CFG181;
  input CFG208;
  input CFG211;
  input CFG178;
  input CBE_I5;
  input CFG212;
  input CFG182;
  input CFG209;
  input CFG179;
  input CBE_I6;
  input CFG213;
  input CFG183;
  input CBE_I7;
  input CFG214;
  input CFG184;
  input CFG185;
  input CFG215;
  input CFG186;
  input CFG216;
  input CFG190;
  input CFG220;
  input CFG217;
  input CFG187;
  input CFG191;
  input CFG221;
  input CFG218;
  input CFG188;
  input CFG192;
  input CFG222;
  input CFG219;
  input CFG189;
  input CFG193;
  input CFG223;
  input CFG194;
  input CFG224;
  input CFG195;
  input CFG225;
  input CFG196;
  input CFG226;
  input CFG197;
  input CFG230;
  input CFG227;
  input CFG198;
  input CFG231;
  input CFG228;
  input CFG199;
  input CFG232;
  input CFG229;
  input CFG233;
  output B_BUSY;
  input CFG234;
  input CFG235;
  input CFG236;
  input CFG237;
  input CFG240;
  input CFG238;
  output CFG_VLD;
  input CFG241;
  input CFG239;
  input CFG242;
  input CFG243;
  output M_DATA;
  input CFG244;
  input CFG245;
  input CFG246;
  input CFG247;
  input CFG250;
  input CFG248;
  input CFG251;
  input CFG249;
  input CFG252;
  input CFG253;
  output IRDYQ_N;
  input CFG254;
  input CFG255;
  input SERR_I;
  output CBE_O0;
  output OE_PAR;
  output CBE_O1;
  output CBE_O2;
  input REQUEST;
  output CBE_O3;
  output CBE_O4;
  output CBE_O5;
  output CBE_O6;
  output CBE_O7;
  output OE_ADO_LB64;
  output OE_REQ64;
  input KEEPOUT;
  output OE_INTA;
  input REQUESTHOLD;
  input S_ABORT;
  output ADDR0;
  output OE_PAR64;
  output ADDR1;
  output ADDR2;
  output ADDR3;
  output ADDR4;
  output ADDR5;
  output ADDR6;
  output BACKOFF;
  output ADDR7;
  output ADDR8;
  output OE_ADO_T64;
  output ADDR9;
  output CFG_HIT;
  output OE_TRDY;
  input SUB_DATA0;
  input SUB_DATA1;
  input SUB_DATA2;
  input SUB_DATA3;
  input SUB_DATA4;
  input SUB_DATA5;
  input SUB_DATA6;
  output OE_CBE64;
  input SUB_DATA7;
  input SUB_DATA8;
  input SUB_DATA9;
  output FRAMEQ_N;
  output OE_ADO_LB;
  output S_DATA;
  output OE_ADO_LT;
// synthesis translate_off
  wire \$1N4834 ;
  wire \$5N3772 ;
  wire \$5N3783 ;
  wire \$6N1151 ;
  wire \$6N1152 ;
  wire \$6N1153 ;
  wire \$6N1154 ;
  wire \$6N1155 ;
  wire \$6N1156 ;
  wire \$6N1173 ;
  wire \$7N143 ;
  wire \$7N147 ;
  wire \$7N148 ;
  wire \$7N149 ;
  wire \$7N152 ;
  wire \$7N156 ;
  wire \$7N160 ;
  wire \$7N163 ;
  wire \$7N583 ;
  wire \$7N621 ;
  wire \$7N625 ;
  wire \$7N745 ;
  wire \$7N855 ;
  wire \$7N859 ;
  wire \0BR0 ;
  wire \0BR1 ;
  wire \0BR10 ;
  wire \0BR11 ;
  wire \0BR12 ;
  wire \0BR13 ;
  wire \0BR14 ;
  wire \0BR15 ;
  wire \0BR16 ;
  wire \0BR17 ;
  wire \0BR18 ;
  wire \0BR19 ;
  wire \0BR2 ;
  wire \0BR20 ;
  wire \0BR21 ;
  wire \0BR22 ;
  wire \0BR23 ;
  wire \0BR24 ;
  wire \0BR25 ;
  wire \0BR26 ;
  wire \0BR27 ;
  wire \0BR28 ;
  wire \0BR29 ;
  wire \0BR3 ;
  wire \0BR30 ;
  wire \0BR31 ;
  wire \0BR4 ;
  wire \0BR5 ;
  wire \0BR6 ;
  wire \0BR7 ;
  wire \0BR8 ;
  wire \0BR9 ;
  wire \1BR0 ;
  wire \1BR1 ;
  wire \1BR10 ;
  wire \1BR11 ;
  wire \1BR12 ;
  wire \1BR13 ;
  wire \1BR14 ;
  wire \1BR15 ;
  wire \1BR16 ;
  wire \1BR17 ;
  wire \1BR18 ;
  wire \1BR19 ;
  wire \1BR2 ;
  wire \1BR20 ;
  wire \1BR21 ;
  wire \1BR22 ;
  wire \1BR23 ;
  wire \1BR24 ;
  wire \1BR25 ;
  wire \1BR26 ;
  wire \1BR27 ;
  wire \1BR28 ;
  wire \1BR29 ;
  wire \1BR3 ;
  wire \1BR30 ;
  wire \1BR31 ;
  wire \1BR4 ;
  wire \1BR5 ;
  wire \1BR6 ;
  wire \1BR7 ;
  wire \1BR8 ;
  wire \1BR9 ;
  wire \2BR0 ;
  wire \2BR1 ;
  wire \2BR10 ;
  wire \2BR11 ;
  wire \2BR12 ;
  wire \2BR13 ;
  wire \2BR14 ;
  wire \2BR15 ;
  wire \2BR16 ;
  wire \2BR17 ;
  wire \2BR18 ;
  wire \2BR19 ;
  wire \2BR2 ;
  wire \2BR20 ;
  wire \2BR21 ;
  wire \2BR22 ;
  wire \2BR23 ;
  wire \2BR24 ;
  wire \2BR25 ;
  wire \2BR26 ;
  wire \2BR27 ;
  wire \2BR28 ;
  wire \2BR29 ;
  wire \2BR3 ;
  wire \2BR30 ;
  wire \2BR31 ;
  wire \2BR4 ;
  wire \2BR5 ;
  wire \2BR6 ;
  wire \2BR7 ;
  wire \2BR8 ;
  wire \2BR9 ;
  wire \ACK64- ;
  wire ACK64_CE;
  wire NlwRenamedSig_OI_ADDR0;
  wire NlwRenamedSig_OI_ADDR1;
  wire NlwRenamedSig_OI_ADDR10;
  wire NlwRenamedSig_OI_ADDR11;
  wire NlwRenamedSig_OI_ADDR12;
  wire NlwRenamedSig_OI_ADDR13;
  wire NlwRenamedSig_OI_ADDR14;
  wire NlwRenamedSig_OI_ADDR15;
  wire NlwRenamedSig_OI_ADDR16;
  wire NlwRenamedSig_OI_ADDR17;
  wire NlwRenamedSig_OI_ADDR18;
  wire NlwRenamedSig_OI_ADDR19;
  wire NlwRenamedSig_OI_ADDR2;
  wire NlwRenamedSig_OI_ADDR20;
  wire NlwRenamedSig_OI_ADDR21;
  wire NlwRenamedSig_OI_ADDR22;
  wire NlwRenamedSig_OI_ADDR23;
  wire NlwRenamedSig_OI_ADDR24;
  wire NlwRenamedSig_OI_ADDR25;
  wire NlwRenamedSig_OI_ADDR26;
  wire NlwRenamedSig_OI_ADDR27;
  wire NlwRenamedSig_OI_ADDR28;
  wire NlwRenamedSig_OI_ADDR29;
  wire NlwRenamedSig_OI_ADDR3;
  wire NlwRenamedSig_OI_ADDR30;
  wire NlwRenamedSig_OI_ADDR31;
  wire NlwRenamedSig_OI_ADDR4;
  wire NlwRenamedSig_OI_ADDR5;
  wire NlwRenamedSig_OI_ADDR6;
  wire NlwRenamedSig_OI_ADDR7;
  wire NlwRenamedSig_OI_ADDR8;
  wire NlwRenamedSig_OI_ADDR9;
  wire ADDR_BE;
  wire NlwRenamedSig_OI_ADDR_VLD;
  wire ADDR_VLD0;
  wire ADDR_VLD1;
  wire ADDR_VLD64;
  wire ADOUT0;
  wire ADOUT1;
  wire ADOUT10;
  wire ADOUT11;
  wire ADOUT12;
  wire ADOUT13;
  wire ADOUT14;
  wire ADOUT15;
  wire ADOUT16;
  wire ADOUT17;
  wire ADOUT18;
  wire ADOUT19;
  wire ADOUT2;
  wire ADOUT20;
  wire ADOUT21;
  wire ADOUT22;
  wire ADOUT23;
  wire ADOUT24;
  wire ADOUT25;
  wire ADOUT26;
  wire ADOUT27;
  wire ADOUT28;
  wire ADOUT29;
  wire ADOUT3;
  wire ADOUT30;
  wire ADOUT31;
  wire ADOUT32;
  wire ADOUT33;
  wire ADOUT34;
  wire ADOUT35;
  wire ADOUT36;
  wire ADOUT37;
  wire ADOUT38;
  wire ADOUT39;
  wire ADOUT4;
  wire ADOUT40;
  wire ADOUT41;
  wire ADOUT42;
  wire ADOUT43;
  wire ADOUT44;
  wire ADOUT45;
  wire ADOUT46;
  wire ADOUT47;
  wire ADOUT48;
  wire ADOUT49;
  wire ADOUT5;
  wire ADOUT50;
  wire ADOUT51;
  wire ADOUT52;
  wire ADOUT53;
  wire ADOUT54;
  wire ADOUT55;
  wire ADOUT56;
  wire ADOUT57;
  wire ADOUT58;
  wire ADOUT59;
  wire ADOUT6;
  wire ADOUT60;
  wire ADOUT61;
  wire ADOUT62;
  wire ADOUT63;
  wire ADOUT7;
  wire ADOUT8;
  wire ADOUT9;
  wire APERR_N;
  wire ATTEMPT64;
  wire BACKOFF_INT;
  wire BAR0_T;
  wire BAR1_T;
  wire BAR2_T;
  wire BAR3;
  wire BAR4;
  wire BAR5;
  wire BAR6;
  wire BAR7;
  wire NlwRenamedSig_OI_BASE_HIT0;
  wire NlwRenamedSig_OI_BASE_HIT1;
  wire NlwRenamedSig_OI_BASE_HIT2;
  wire BASE_HIT2_INT;
  wire NlwRenamedSig_OI_BASE_HIT3;
  wire NlwRenamedSig_OI_BASE_HIT4;
  wire NlwRenamedSig_OI_BASE_HIT5;
  wire NlwRenamedSig_OI_BASE_HIT6;
  wire NlwRenamedSig_OI_BASE_HIT7;
  wire BH64_0;
  wire BH64_1;
  wire BH64_2;
  wire BH64_2_INT;
  wire B_BUSY_INT;
  wire CBEOUT0;
  wire CBEOUT1;
  wire CBEOUT2;
  wire CBEOUT3;
  wire CBEOUT4;
  wire CBEOUT5;
  wire CBEOUT6;
  wire CBEOUT7;
  wire CE0_0;
  wire CE0_1;
  wire CE0_2;
  wire CE0_3;
  wire CE10_0;
  wire CE10_1;
  wire CE10_2;
  wire CE10_3;
  wire CE11_0;
  wire CE11_1;
  wire CE11_2;
  wire CE11_3;
  wire CE12_0;
  wire CE12_1;
  wire CE12_2;
  wire CE12_3;
  wire CE13_0;
  wire CE13_1;
  wire CE13_2;
  wire CE13_3;
  wire CE14_0;
  wire CE14_1;
  wire CE14_2;
  wire CE14_3;
  wire CE15_0;
  wire CE15_1;
  wire CE15_2;
  wire CE15_3;
  wire CE1_0;
  wire CE1_1;
  wire CE1_2;
  wire CE1_3;
  wire CE2_0;
  wire CE2_1;
  wire CE2_2;
  wire CE2_3;
  wire CE3_0;
  wire CE3_1;
  wire CE3_2;
  wire CE3_3;
  wire CE4_0;
  wire CE4_1;
  wire CE4_2;
  wire CE4_3;
  wire CE5_0;
  wire CE5_1;
  wire CE5_2;
  wire CE5_3;
  wire CE6_0;
  wire CE6_1;
  wire CE6_2;
  wire CE6_3;
  wire CE7_0;
  wire CE7_1;
  wire CE7_2;
  wire CE7_3;
  wire CE8_0;
  wire CE8_1;
  wire CE8_2;
  wire CE8_3;
  wire CE9_0;
  wire CE9_1;
  wire CE9_2;
  wire CE9_3;
  wire NlwRenamedSig_OI_CFG_HIT;
  wire NlwRenamedSig_OI_CFG_VLD;
  wire NlwRenamedSig_OI_CSR0;
  wire NlwRenamedSig_OI_CSR1;
  wire NlwRenamedSig_OI_CSR10;
  wire NlwRenamedSig_OI_CSR11;
  wire NlwRenamedSig_OI_CSR12;
  wire NlwRenamedSig_OI_CSR13;
  wire NlwRenamedSig_OI_CSR14;
  wire NlwRenamedSig_OI_CSR15;
  wire NlwRenamedSig_OI_CSR16;
  wire NlwRenamedSig_OI_CSR17;
  wire NlwRenamedSig_OI_CSR18;
  wire NlwRenamedSig_OI_CSR19;
  wire NlwRenamedSig_OI_CSR2;
  wire NlwRenamedSig_OI_CSR20;
  wire NlwRenamedSig_OI_CSR21;
  wire NlwRenamedSig_OI_CSR22;
  wire NlwRenamedSig_OI_CSR23;
  wire NlwRenamedSig_OI_CSR24;
  wire NlwRenamedSig_OI_CSR25;
  wire NlwRenamedSig_OI_CSR26;
  wire NlwRenamedSig_OI_CSR27;
  wire NlwRenamedSig_OI_CSR28;
  wire NlwRenamedSig_OI_CSR29;
  wire NlwRenamedSig_OI_CSR3;
  wire NlwRenamedSig_OI_CSR30;
  wire NlwRenamedSig_OI_CSR31;
  wire NlwRenamedSig_OI_CSR32;
  wire NlwRenamedSig_OI_CSR33;
  wire NlwRenamedSig_OI_CSR34;
  wire NlwRenamedSig_OI_CSR35;
  wire NlwRenamedSig_OI_CSR36;
  wire NlwRenamedSig_OI_CSR37;
  wire NlwRenamedSig_OI_CSR38;
  wire NlwRenamedSig_OI_CSR39;
  wire NlwRenamedSig_OI_CSR4;
  wire NlwRenamedSig_OI_CSR5;
  wire NlwRenamedSig_OI_CSR6;
  wire NlwRenamedSig_OI_CSR7;
  wire NlwRenamedSig_OI_CSR8;
  wire NlwRenamedSig_OI_CSR9;
  wire \DEVSEL- ;
  wire DEVSEL_CE;
  wire DP64_T;
  wire DR_BUS_INT;
  wire EOT;
  wire EX;
  wire FAIL64_INT;
  wire FAIL_ADH32;
  wire FAIL_ADH33;
  wire FAIL_ADH34;
  wire FAIL_ADH35;
  wire FAIL_ADH36;
  wire FAIL_ADH37;
  wire FAIL_ADH38;
  wire FAIL_ADH39;
  wire FAIL_ADH40;
  wire FAIL_ADH41;
  wire FAIL_ADH42;
  wire FAIL_ADH43;
  wire FAIL_ADH44;
  wire FAIL_ADH45;
  wire FAIL_ADH46;
  wire FAIL_ADH47;
  wire FAIL_ADH48;
  wire FAIL_ADH49;
  wire FAIL_ADH50;
  wire FAIL_ADH51;
  wire FAIL_ADH52;
  wire FAIL_ADH53;
  wire FAIL_ADH54;
  wire FAIL_ADH55;
  wire FAIL_ADH56;
  wire FAIL_ADH57;
  wire FAIL_ADH58;
  wire FAIL_ADH59;
  wire FAIL_ADH60;
  wire FAIL_ADH61;
  wire FAIL_ADH62;
  wire FAIL_ADH63;
  wire FAIL_CBH4;
  wire FAIL_CBH5;
  wire FAIL_CBH6;
  wire FAIL_CBH7;
  wire FAKE_GTS_13003;
  wire \FRAME- ;
  wire FRAME_CE;
  wire \GNT- ;
  wire HAS_IO;
  wire HAS_MEM;
  wire IDLE_DUP;
  wire IDLE_INT;
  wire IDSEL;
  wire IDSEL_O;
  wire \IFRAME_I- ;
  wire \IIRDY_I- ;
  wire INTACK;
  wire INTACKQ;
  wire IPWIN;
  wire IPWIN64;
  wire \IRDY- ;
  wire IRDY_CE;
  wire IRDY_F;
  wire IRDY_M;
  wire IREG0;
  wire IREG1;
  wire IREG10;
  wire IREG11;
  wire IREG12;
  wire IREG13;
  wire IREG14;
  wire IREG15;
  wire IREG16;
  wire IREG17;
  wire IREG18;
  wire IREG19;
  wire IREG2;
  wire IREG20;
  wire IREG21;
  wire IREG22;
  wire IREG23;
  wire IREG24;
  wire IREG25;
  wire IREG26;
  wire IREG27;
  wire IREG28;
  wire IREG29;
  wire IREG3;
  wire IREG30;
  wire IREG31;
  wire IREG4;
  wire IREG5;
  wire IREG6;
  wire IREG7;
  wire IREG8;
  wire IREG9;
  wire \IREQ64_I- ;
  wire I_IDLE_INT;
  wire MD0;
  wire MD1;
  wire MD10;
  wire MD11;
  wire MD12;
  wire MD13;
  wire MD14;
  wire MD15;
  wire MD16;
  wire MD17;
  wire MD18;
  wire MD19;
  wire MD2;
  wire MD20;
  wire MD21;
  wire MD22;
  wire MD23;
  wire MD24;
  wire MD25;
  wire MD26;
  wire MD27;
  wire MD28;
  wire MD29;
  wire MD3;
  wire MD30;
  wire MD31;
  wire MD4;
  wire MD5;
  wire MD6;
  wire MD7;
  wire MD8;
  wire MD9;
  wire MIKELOVEJOY;
  wire M_CBE_INT0;
  wire M_CBE_INT1;
  wire M_CBE_INT2;
  wire M_CBE_INT3;
  wire M_CBE_INT4;
  wire M_CBE_INT5;
  wire M_CBE_INT6;
  wire M_CBE_INT7;
  wire M_DATA_INT;
  wire M_ENABLE;
  wire M_FIRST;
  wire NlwRenamedSig_OI_M_SRC_EN;
  wire NEWDATA;
  wire NL3;
  wire NL4;
  wire NL5;
  wire NL6;
  wire NL7;
  wire NL_MEM0;
  wire NL_MEM1;
  wire NL_MEM2;
  wire NL_MEM3;
  wire NL_MEM4;
  wire NL_MEM5;
  wire NL_MEM6;
  wire NL_MEM7;
  wire \NS_ACK64- ;
  wire NS_BASE_HIT0;
  wire NS_BASE_HIT1;
  wire NS_BASE_HIT2;
  wire NS_BASE_HIT2_INT;
  wire NS_BH64_0;
  wire NS_BH64_1;
  wire NS_BH64_2;
  wire NS_BH64_2_INT;
  wire \NS_DEVSEL- ;
  wire \NS_FRAME- ;
  wire NS_IDSEL;
  wire \NS_IRDY- ;
  wire NS_OE_PERR_T;
  wire NS_PAR;
  wire NS_PAR64;
  wire \NS_PERR- ;
  wire \NS_REQ64- ;
  wire \NS_SERR- ;
  wire \NS_STOP- ;
  wire \NS_TRDY- ;
  wire OE0;
  wire OE1;
  wire OE10;
  wire OE11;
  wire OE12;
  wire OE13;
  wire OE14;
  wire OE15;
  wire OE2;
  wire OE3;
  wire OE4;
  wire OE5;
  wire OE6;
  wire OE7;
  wire OE8;
  wire OE9;
  wire OE_ADI;
  wire OE_ADI64;
  wire NlwRenamedSig_OI_OE_ADO_B;
  wire NlwRenamedSig_OI_OE_ADO_B64;
  wire NlwRenamedSig_OI_OE_ADO_LB;
  wire NlwRenamedSig_OI_OE_ADO_LB64;
  wire NlwRenamedSig_OI_OE_ADO_LT;
  wire NlwRenamedSig_OI_OE_ADO_LT64;
  wire NlwRenamedSig_OI_OE_ADO_T;
  wire NlwRenamedSig_OI_OE_ADO_T64;
  wire OE_AD_T_B;
  wire OE_AD_T_B64;
  wire OE_AD_T_LB;
  wire OE_AD_T_LB64;
  wire OE_AD_T_LT;
  wire OE_AD_T_LT64;
  wire OE_AD_T_T;
  wire OE_AD_T_T64;
  wire NlwRenamedSig_OI_OE_CBE;
  wire NlwRenamedSig_OI_OE_CBE64;
  wire NlwRenamedSig_OI_OE_PAR;
  wire NlwRenamedSig_OI_OE_PAR64;
  wire OE_ROM;
  wire OLDKEEPOUT;
  wire OUT_SEL;
  wire OUT_SEL64;
  wire PAR_CE;
  wire PCI_CE;
  wire NlwRenamedSig_OI_PCI_CMD0;
  wire NlwRenamedSig_OI_PCI_CMD1;
  wire NlwRenamedSig_OI_PCI_CMD10;
  wire NlwRenamedSig_OI_PCI_CMD11;
  wire NlwRenamedSig_OI_PCI_CMD12;
  wire NlwRenamedSig_OI_PCI_CMD13;
  wire NlwRenamedSig_OI_PCI_CMD14;
  wire NlwRenamedSig_OI_PCI_CMD15;
  wire NlwRenamedSig_OI_PCI_CMD2;
  wire NlwRenamedSig_OI_PCI_CMD3;
  wire NlwRenamedSig_OI_PCI_CMD4;
  wire NlwRenamedSig_OI_PCI_CMD5;
  wire NlwRenamedSig_OI_PCI_CMD6;
  wire NlwRenamedSig_OI_PCI_CMD7;
  wire NlwRenamedSig_OI_PCI_CMD8;
  wire NlwRenamedSig_OI_PCI_CMD9;
  wire \PERR- ;
  wire PERR_EN;
  wire \REQ64- ;
  wire REQ64_CE;
  wire NlwRenamedSig_OI_RST;
  wire \SERR- ;
  wire SERR_EN;
  wire SERR_O;
  wire SET0;
  wire SET1;
  wire SET10;
  wire SET11;
  wire SET12;
  wire SET13;
  wire SET14;
  wire SET15;
  wire SET2;
  wire SET3;
  wire SET4;
  wire SET5;
  wire SET6;
  wire SET7;
  wire SET8;
  wire SET9;
  wire SHADOW0;
  wire SHADOW1;
  wire SHADOW10;
  wire SHADOW11;
  wire SHADOW12;
  wire SHADOW13;
  wire SHADOW14;
  wire SHADOW15;
  wire SHADOW16;
  wire SHADOW17;
  wire SHADOW18;
  wire SHADOW19;
  wire SHADOW2;
  wire SHADOW20;
  wire SHADOW21;
  wire SHADOW22;
  wire SHADOW23;
  wire SHADOW24;
  wire SHADOW25;
  wire SHADOW26;
  wire SHADOW27;
  wire SHADOW28;
  wire SHADOW29;
  wire SHADOW3;
  wire SHADOW30;
  wire SHADOW31;
  wire SHADOW32;
  wire SHADOW33;
  wire SHADOW34;
  wire SHADOW35;
  wire SHADOW36;
  wire SHADOW37;
  wire SHADOW38;
  wire SHADOW39;
  wire SHADOW4;
  wire SHADOW40;
  wire SHADOW41;
  wire SHADOW42;
  wire SHADOW43;
  wire SHADOW44;
  wire SHADOW45;
  wire SHADOW46;
  wire SHADOW47;
  wire SHADOW48;
  wire SHADOW49;
  wire SHADOW5;
  wire SHADOW50;
  wire SHADOW51;
  wire SHADOW52;
  wire SHADOW53;
  wire SHADOW54;
  wire SHADOW55;
  wire SHADOW56;
  wire SHADOW57;
  wire SHADOW58;
  wire SHADOW59;
  wire SHADOW6;
  wire SHADOW60;
  wire SHADOW61;
  wire SHADOW62;
  wire SHADOW63;
  wire SHADOW7;
  wire SHADOW8;
  wire SHADOW9;
  wire SHADOW_CBE0;
  wire SHADOW_CBE1;
  wire SHADOW_CBE2;
  wire SHADOW_CBE3;
  wire SHADOW_CBE4;
  wire SHADOW_CBE5;
  wire SHADOW_CBE6;
  wire SHADOW_CBE7;
  wire SHADOW_CE;
  wire SHADOW_CE64;
  wire \STOP- ;
  wire STOP_CE;
  wire NlwRenamedSig_OI_S_CBE0;
  wire NlwRenamedSig_OI_S_CBE1;
  wire NlwRenamedSig_OI_S_CBE2;
  wire NlwRenamedSig_OI_S_CBE3;
  wire NlwRenamedSig_OI_S_CBE4;
  wire NlwRenamedSig_OI_S_CBE5;
  wire NlwRenamedSig_OI_S_CBE6;
  wire NlwRenamedSig_OI_S_CBE7;
  wire S_CYCLE64_INT;
  wire S_DATA_INT;
  wire S_FIRST;
  wire NlwRenamedSig_OI_S_WRDN;
  wire S_WRDN_DUP;
  wire \TACK64_I- ;
  wire \TDEVSEL_I- ;
  wire NlwRenamedSig_OI_TIME_OUT;
  wire TPWIN;
  wire TPWIN64;
  wire \TRDY- ;
  wire TRDY_CE;
  wire TRDY_F;
  wire TRDY_M;
  wire \TSTOP_I- ;
  wire \TTRDY_I- ;
  wire TURN_AR_INT;
  wire \MASTER/$4N3252 ;
  wire \MASTER/REG_0CH26 ;
  wire \MASTER/REG_0CH25 ;
  wire \MASTER/REG_0CH24 ;
  wire \MASTER/REG_0CH23 ;
  wire \MASTER/REG_0CH22 ;
  wire \MASTER/REG_0CH19 ;
  wire \MASTER/REG_0CH21 ;
  wire \MASTER/REG_0CH18 ;
  wire \MASTER/REG_0CH20 ;
  wire \MASTER/REG_0CH17 ;
  wire \MASTER/REG_0CH16 ;
  wire \MASTER/REG_0CH7 ;
  wire \MASTER/REG_0CH6 ;
  wire \MASTER/REG_0CH5 ;
  wire \MASTER/REG_0CH4 ;
  wire \MASTER/REG_0CH3 ;
  wire \MASTER/REG_0CH2 ;
  wire \MASTER/REG_0CH1 ;
  wire \MASTER/REG_0CH0 ;
  wire \MASTER/REG_0CH29 ;
  wire \MASTER/REG_0CH31 ;
  wire \MASTER/REG_0CH28 ;
  wire \MASTER/REG_0CH30 ;
  wire \MASTER/REG_0CH27 ;
  wire \MASTER/REG_0CH8 ;
  wire \MASTER/REG_0CH9 ;
  wire \MASTER/REG_0CH10 ;
  wire \MASTER/REG_0CH11 ;
  wire \MASTER/REG_0CH12 ;
  wire \MASTER/REG_0CH13 ;
  wire \MASTER/REG_0CH14 ;
  wire \MASTER/REG_0CH15 ;
  wire \MASTER/LAT_TIME7 ;
  wire \MASTER/LAT_TIME6 ;
  wire \MASTER/LAT_TIME5 ;
  wire \MASTER/LAT_TIME4 ;
  wire \MASTER/LAT_TIME3 ;
  wire \MASTER/LAT_TIME2 ;
  wire \MASTER/LAT_TIME1 ;
  wire \MASTER/LAT_TIME0 ;
  wire \MASTER/CNT_VAL7 ;
  wire \MASTER/CNT_VAL6 ;
  wire \MASTER/CNT_VAL5 ;
  wire \MASTER/CNT_VAL4 ;
  wire \MASTER/CNT_VAL3 ;
  wire \MASTER/CNT_VAL2 ;
  wire \MASTER/CNT_VAL1 ;
  wire \MASTER/CNT_VAL0 ;
  wire \MASTER/$4N3302 ;
  wire \MASTER/REQ- ;
  wire \MASTER/NS_GNT- ;
  wire \MASTER/GNT_O ;
  wire \MASTER/NS_IREAD64 ;
  wire \MASTER/IREAD64 ;
  wire \MASTER/$4N3030 ;
  wire \MASTER/$4N3021 ;
  wire \MASTER/IREQ64- ;
  wire \MASTER/IREQ_I- ;
  wire \MASTER/NS_REQ- ;
  wire \MASTER/IREQ- ;
  wire \MASTER/S_TAR ;
  wire \MASTER/IIRDY- ;
  wire \MASTER/REQUEST64 ;
  wire \MASTER/REQUEST ;
  wire \MASTER/M_ENABLE ;
  wire \MASTER/DEV_TO ;
  wire \MASTER/IFRAME- ;
  wire \MASTER/I_IDLE/VALIDREQ ;
  wire \MASTER/I_IDLE/ADDR_GNT ;
  wire \MASTER/I_IDLE/$1N2776 ;
  wire \MASTER/I_IDLE/EQ-C ;
  wire \MASTER/I_IDLE/EQ-B ;
  wire \MASTER/I_IDLE/PRE_C2 ;
  wire \MASTER/I_IDLE/EQ-A ;
  wire \MASTER/I_IDLE/M_DATA_C1 ;
  wire \MASTER/I_IDLE/M_DATA_C2 ;
  wire \MASTER/I_IDLE/M_DATA_AND_DR_BUS ;
  wire \MASTER/I_IDLE/I_IDLE_ADDR_GNT ;
  wire \MASTER/I_IDLE/NS_I_IDLE ;
  wire \MASTER/ADDR/$1N2628 ;
  wire \MASTER/ADDR/NS_MAN ;
  wire \MASTER/ADDR/$1N2603 ;
  wire \MASTER/ADDR/M_ADDR_DEAD ;
  wire \MASTER/ADDR/NS_ABE ;
  wire \MASTER/DR_BUS/$1N2925 ;
  wire \MASTER/DR_BUS/BBBRGH ;
  wire \MASTER/DR_BUS/$1N2812 ;
  wire \MASTER/DR_BUS/$1N2820 ;
  wire \MASTER/DR_BUS/AAARGH ;
  wire \MASTER/DR_BUS/$1N2745 ;
  wire \MASTER/DR_BUS/$1N2793 ;
  wire \MASTER/DR_BUS/COMMON-B ;
  wire \MASTER/DR_BUS/COMMON-A ;
  wire \MASTER/DR_BUS/COND ;
  wire \MASTER/DR_BUS/EQN-B0 ;
  wire \MASTER/DR_BUS/$1N2718 ;
  wire \MASTER/DR_BUS/$1N2720 ;
  wire \MASTER/DR_BUS/EQN-A0 ;
  wire \MASTER/DR_BUS/$1N2700 ;
  wire \MASTER/DR_BUS/EQN-A1 ;
  wire \MASTER/DR_BUS/EQN-B1 ;
  wire \MASTER/DR_BUS/NS_1 ;
  wire \MASTER/DR_BUS/NS_0 ;
  wire \MASTER/DR_BUS/NS_DR_BUS ;
  wire \MASTER/DR_BUS/$1I2908/M1 ;
  wire \MASTER/DR_BUS/$1I2908/M0 ;
  wire \MASTER/DR_BUS/$1I2917/M1 ;
  wire \MASTER/DR_BUS/$1I2917/M0 ;
  wire \MASTER/DR_BUS/$1I2927/$1N2216 ;
  wire \MASTER/M_DATA/$1N2519 ;
  wire \MASTER/M_DATA/EQN-A ;
  wire \MASTER/M_DATA/EQN_B ;
  wire \MASTER/M_DATA/$1N2507 ;
  wire \MASTER/M_DATA/NS_MDATA ;
  wire \MASTER/$1I2914/END_OF_XFER ;
  wire \MASTER/$1I2914/$1N2929 ;
  wire \MASTER/$1I2914/$1N2938 ;
  wire \MASTER/$1I2914/$1N2959 ;
  wire \MASTER/$1I2914/M_DATA_Q ;
  wire \MASTER/$1I2914/REQUEST64Q ;
  wire \MASTER/$1I2914/$1N2897 ;
  wire \MASTER/$1I2914/LOCKOUT ;
  wire \MASTER/$1I2914/$1N2884 ;
  wire \MASTER/$1I2914/SCG32 ;
  wire \MASTER/$1I2914/SCG64 ;
  wire \MASTER/$1I2914/$1N2894 ;
  wire \MASTER/$1I2914/ADDR_BE_Q ;
  wire \MASTER/$1I2914/$1N2881 ;
  wire \MASTER/$1I2914/CANCEL ;
  wire \MASTER/$1I2914/$1I2853/$1N2215 ;
  wire \MASTER/$1I2914/$1I2853/D ;
  wire \MASTER/$1I2914/$1I2864/$1N2215 ;
  wire \MASTER/$1I2914/$1I2864/D ;
  wire \MASTER/$1I2914/$1I2932/$1N2215 ;
  wire \MASTER/$1I2914/$1I2932/D ;
  wire \MASTER/FRAME/$2N3531 ;
  wire \MASTER/FRAME/DTO ;
  wire \MASTER/FRAME/$2N3521 ;
  wire \MASTER/FRAME/$2N3475 ;
  wire \MASTER/FRAME/$2N3449 ;
  wire \MASTER/FRAME/$2N3450 ;
  wire \MASTER/FRAME/DONE_1 ;
  wire \MASTER/FRAME/INITIAL ;
  wire \MASTER/FRAME/DONE_0 ;
  wire \MASTER/FRAME/$1N3468 ;
  wire \MASTER/FRAME/$1N3369 ;
  wire \MASTER/FRAME/IRDY_64 ;
  wire \MASTER/FRAME/NS_S_1 ;
  wire \MASTER/FRAME/KO_T_0 ;
  wire \MASTER/FRAME/KO_T_1 ;
  wire \MASTER/FRAME/NS_S_0 ;
  wire \MASTER/FRAME/TURN_ON ;
  wire \MASTER/FRAME/FEEDBACK ;
  wire \MASTER/FRAME/$1I3467/M1 ;
  wire \MASTER/FRAME/$1I3467/M0 ;
  wire \MASTER/FRAME/$2I3559/M1 ;
  wire \MASTER/FRAME/$2I3559/M0 ;
  wire \MASTER/IRDY/EQN-F ;
  wire \MASTER/IRDY/$2N3385 ;
  wire \MASTER/IRDY/M_FIRSTIN ;
  wire \MASTER/IRDY/$2N3355 ;
  wire \MASTER/IRDY/$2N3294 ;
  wire \MASTER/IRDY/M_FIRST1 ;
  wire \MASTER/IRDY/M_FIRST0 ;
  wire \MASTER/IRDY/$2N3383 ;
  wire \MASTER/IRDY/END_OF_INIT ;
  wire \MASTER/IRDY/M_DATA_Q ;
  wire \MASTER/IRDY/$1N3756 ;
  wire \MASTER/IRDY/EQN-G ;
  wire \MASTER/IRDY/$1N3772 ;
  wire \MASTER/IRDY/$1N3721 ;
  wire \MASTER/IRDY/$1N3502 ;
  wire \MASTER/IRDY/WS_A_1 ;
  wire \MASTER/IRDY/WS_A_0 ;
  wire \MASTER/IRDY/$1N3493 ;
  wire \MASTER/IRDY/NS_1 ;
  wire \MASTER/IRDY/ALLOWED ;
  wire \MASTER/IRDY/CORE_READY ;
  wire \MASTER/IRDY/NS_0 ;
  wire \MASTER/IRDY/EQN-E ;
  wire \MASTER/IRDY/$1I3227/M1 ;
  wire \MASTER/IRDY/$1I3227/M0 ;
  wire \MASTER/IRDY/$1I3492/M1 ;
  wire \MASTER/IRDY/$1I3492/M0 ;
  wire \MASTER/IRDY/$1I3563/$1N2216 ;
  wire \MASTER/IRDY/$2I3285/M1 ;
  wire \MASTER/IRDY/$2I3285/M0 ;
  wire \MASTER/REQ/EXT ;
  wire \MASTER/REQ/S_TAR_OR ;
  wire \MASTER/REQ/NORM1 ;
  wire \MASTER/REQ/NORM2 ;
  wire \MASTER/REQ/SOXFER ;
  wire \MASTER/REQ/REQ_BUS ;
  wire \MASTER/REQ/$1N2737 ;
  wire \MASTER/REQ/M_DATA_Q ;
  wire \MASTER/REQ/X ;
  wire \MASTER/REQ/S_TARQ ;
  wire \MASTER/REQ/Y ;
  wire \MASTER/REQ/$1I2708/$1N2215 ;
  wire \MASTER/REQ/$1I2708/D ;
  wire \MASTER/REQ64/DONE_0 ;
  wire \MASTER/REQ64/$2N3399 ;
  wire \MASTER/REQ64/INITIAL ;
  wire \MASTER/REQ64/$2N3428 ;
  wire \MASTER/REQ64/$2N3430 ;
  wire \MASTER/REQ64/$2N3429 ;
  wire \MASTER/REQ64/DTO ;
  wire \MASTER/REQ64/DONE_1 ;
  wire \MASTER/REQ64/$2N3396 ;
  wire \MASTER/REQ64/FEEDBACK ;
  wire \MASTER/REQ64/$1N3605 ;
  wire \MASTER/REQ64/NS_S_0 ;
  wire \MASTER/REQ64/KO_T_1 ;
  wire \MASTER/REQ64/KO_T_0 ;
  wire \MASTER/REQ64/NS_S_1 ;
  wire \MASTER/REQ64/$1N3615 ;
  wire \MASTER/REQ64/TURN_ON ;
  wire \MASTER/REQ64/IRDY_64 ;
  wire \MASTER/REQ64/$1I3562/M1 ;
  wire \MASTER/REQ64/$1I3562/M0 ;
  wire \MASTER/REQ64/$2I3446/M1 ;
  wire \MASTER/REQ64/$2I3446/M0 ;
  wire \MASTER/XFERFAIL/EQN-X ;
  wire \MASTER/XFERFAIL/SET_FAIL64 ;
  wire \MASTER/XFERFAIL/FEEDBACK ;
  wire \MASTER/XFERFAIL/NS_FAIL64 ;
  wire \MASTER/XFERFAIL/NS_1 ;
  wire \MASTER/XFERFAIL/NS_0 ;
  wire \MASTER/OE_FRAME/$8N4094 ;
  wire \MASTER/OE_FRAME/CE_OER ;
  wire \MASTER/OE_FRAME/NS_OER ;
  wire \MASTER/OE_FRAME/NS_OER_1 ;
  wire \MASTER/OE_FRAME/NS_OER_0 ;
  wire \MASTER/OE_FRAME/$8N4025 ;
  wire \MASTER/OE_FRAME/$8N4024 ;
  wire \MASTER/OE_FRAME/$8N4018 ;
  wire \MASTER/OE_FRAME/$8N4019 ;
  wire \MASTER/OE_FRAME/$8N4080 ;
  wire \MASTER/OE_FRAME/CE_OEF ;
  wire \MASTER/OE_FRAME/$8N3991 ;
  wire \MASTER/OE_FRAME/$8N3986 ;
  wire \MASTER/OE_FRAME/$8N3992 ;
  wire \MASTER/OE_FRAME/$8N3985 ;
  wire \MASTER/OE_FRAME/NS_OEF ;
  wire \MASTER/OE_FRAME/NS_OEF_0 ;
  wire \MASTER/OE_FRAME/NS_OEF_1 ;
  wire \MASTER/OE_FRAME/NS64_1 ;
  wire \MASTER/OE_FRAME/NS64_0 ;
  wire \MASTER/OE_FRAME/$7N3953 ;
  wire \MASTER/OE_FRAME/MISC64_1 ;
  wire \MASTER/OE_FRAME/MISC64_3 ;
  wire \MASTER/OE_FRAME/OE_REQ64_INT_525 ;
  wire \MASTER/OE_FRAME/$7N3948 ;
  wire \MASTER/OE_FRAME/$7N3952 ;
  wire \MASTER/OE_FRAME/$7N3947 ;
  wire \MASTER/OE_FRAME/$7N3949 ;
  wire \MASTER/OE_FRAME/$7N3936 ;
  wire \MASTER/OE_FRAME/$7N3940 ;
  wire \MASTER/OE_FRAME/MISC64_0 ;
  wire \MASTER/OE_FRAME/MISC64_2 ;
  wire \MASTER/OE_FRAME/$7N3955 ;
  wire \MASTER/OE_FRAME/NS64 ;
  wire \MASTER/OE_FRAME/NS_1 ;
  wire \MASTER/OE_FRAME/NS_0 ;
  wire \MASTER/OE_FRAME/$6N3723 ;
  wire \MASTER/OE_FRAME/MISC_1 ;
  wire \MASTER/OE_FRAME/MISC_3 ;
  wire \MASTER/OE_FRAME/OE_FRAME_INT_509 ;
  wire \MASTER/OE_FRAME/$6N3718 ;
  wire \MASTER/OE_FRAME/$6N3722 ;
  wire \MASTER/OE_FRAME/$6N3717 ;
  wire \MASTER/OE_FRAME/$6N3719 ;
  wire \MASTER/OE_FRAME/$6N3707 ;
  wire \MASTER/OE_FRAME/$6N3710 ;
  wire \MASTER/OE_FRAME/MISC_0 ;
  wire \MASTER/OE_FRAME/MISC_2 ;
  wire \MASTER/OE_FRAME/$6N3725 ;
  wire \MASTER/OE_FRAME/NS ;
  wire \MASTER/OE_FRAME/$5N3897 ;
  wire \MASTER/OE_FRAME/$5N3892 ;
  wire \MASTER/OE_FRAME/$5N3876 ;
  wire \MASTER/OE_FRAME/CB64 ;
  wire \MASTER/OE_FRAME/$5N3873 ;
  wire \MASTER/OE_FRAME/$5N3872 ;
  wire \MASTER/OE_FRAME/$5N3871 ;
  wire \MASTER/OE_FRAME/AD_B64 ;
  wire \MASTER/OE_FRAME/AD_LB64 ;
  wire \MASTER/OE_FRAME/$5N3896 ;
  wire \MASTER/OE_FRAME/AD_LT64 ;
  wire \MASTER/OE_FRAME/$5N3895 ;
  wire \MASTER/OE_FRAME/AD_T64 ;
  wire \MASTER/OE_FRAME/$5N3894 ;
  wire \MASTER/OE_FRAME/$5N3874 ;
  wire \MASTER/OE_FRAME/$5N3869 ;
  wire \MASTER/OE_FRAME/$5N3868 ;
  wire \MASTER/OE_FRAME/$5N3870 ;
  wire \MASTER/OE_FRAME/SLOT64 ;
  wire \MASTER/OE_FRAME/CB32 ;
  wire \MASTER/OE_FRAME/AD_B ;
  wire \MASTER/OE_FRAME/$4N3741 ;
  wire \MASTER/OE_FRAME/AD_LB ;
  wire \MASTER/OE_FRAME/$4N3742 ;
  wire \MASTER/OE_FRAME/AD_LT ;
  wire \MASTER/OE_FRAME/$4N3755 ;
  wire \MASTER/OE_FRAME/AD_T ;
  wire \MASTER/OE_FRAME/$4N3754 ;
  wire \MASTER/OE_FRAME/$4N3749 ;
  wire \MASTER/OE_FRAME/$4N3739 ;
  wire \MASTER/OE_FRAME/$4N3738 ;
  wire \MASTER/OE_FRAME/$4N3740 ;
  wire \MASTER/OE_FRAME/SLOT ;
  wire \MASTER/OE_FRAME/EQN-A ;
  wire \MASTER/OE_FRAME/NS_OE_PERR ;
  wire \MASTER/OE_FRAME/SET_OE_PERR ;
  wire \MASTER/OE_FRAME/HOLD_OE_PERR ;
  wire \MASTER/OE_FRAME/START_AD64 ;
  wire \MASTER/OE_FRAME/START_AD ;
  wire \MASTER/OE_FRAME/$1N3716 ;
  wire \MASTER/OE_FRAME/DR_BUS1 ;
  wire \MASTER/OE_FRAME/DUMMY ;
  wire \MASTER/OE_FRAME/DR_BUSQ ;
  wire \MASTER/OE_FRAME/$1N3703 ;
  wire \MASTER/OE_FRAME/REQUEST64Q ;
  wire \MASTER/OE_FRAME/REQUESTQ ;
  wire \MASTER/OE_FRAME/$1N3685 ;
  wire \MASTER/OE_FRAME/$1I3691/$1N2216 ;
  wire \MASTER/OE_FRAME/$1I3717/$1N2216 ;
  wire \MASTER/OE_FRAME/$5I4044/M1 ;
  wire \MASTER/OE_FRAME/$5I4044/M0 ;
  wire \MASTER/OE_FRAME/$5I4045/M1 ;
  wire \MASTER/OE_FRAME/$5I4045/M0 ;
  wire \MASTER/OE_FRAME/$5I4046/M1 ;
  wire \MASTER/OE_FRAME/$5I4046/M0 ;
  wire \MASTER/OE_FRAME/$5I4047/M1 ;
  wire \MASTER/OE_FRAME/$5I4047/M0 ;
  wire \MASTER/OE_FRAME/$5I4048/M1 ;
  wire \MASTER/OE_FRAME/$5I4048/M0 ;
  wire \MASTER/S_TAR/$1N2602 ;
  wire \MASTER/S_TAR/NS_S_TAR ;
  wire \MASTER/DEV_TO/$1N2840 ;
  wire \MASTER/DEV_TO/WAS_SUBTRACTIVE ;
  wire \MASTER/DEV_TO/WAS_NO_RESPONSE ;
  wire \MASTER/DEV_TO/$1N2820 ;
  wire \MASTER/DEV_TO/PASS_TO ;
  wire \MASTER/DEV_TO/WAS_SLOW ;
  wire \MASTER/DEV_TO/WAS_MEDIUM ;
  wire \MASTER/DEV_TO/WAS_FAST ;
  wire \MASTER/DEV_TO/FAST ;
  wire \MASTER/DEV_TO/ADDR ;
  wire \MASTER/DEV_TO/$1I2816/$1N2215 ;
  wire \MASTER/DEV_TO/$1I2816/D ;
  wire \MASTER/DEV_TO/$1I2838/$1N2215 ;
  wire \MASTER/DEV_TO/$1I2838/D ;
  wire \MASTER/$4I3071/$1N2277 ;
  wire \MASTER/$4I3071/$1N2278 ;
  wire \MASTER/$4I3071/$1N2280 ;
  wire \MASTER/GNT_IOB/$1N2286 ;
  wire \MASTER/GNT_IOB/$1N2289 ;
  wire \MASTER/GNT_IOB/$1I2285/$1N2216 ;
  wire \MASTER/GNT_IOB/$1I2288/$1N2216 ;
  wire \MASTER/$4I3148/$1N2216 ;
  wire \MASTER/REQ_IOB/$1N2286 ;
  wire \MASTER/REQ_IOB/$1N2289 ;
  wire \MASTER/REQ_IOB/$1I2285/$1N2216 ;
  wire \MASTER/REQ_IOB/$1I2288/$1N2216 ;
  wire \MASTER/LAT_TIMR/T3 ;
  wire \MASTER/LAT_TIMR/T2 ;
  wire \MASTER/LAT_TIMR/$2N31 ;
  wire \MASTER/LAT_TIMR/$2N13 ;
  wire \MASTER/LAT_TIMR/$1N74 ;
  wire \MASTER/LAT_TIMR/$1N76 ;
  wire \MASTER/LAT_TIMR/TC ;
  wire \MASTER/LAT_TIMR/T000X ;
  wire \MASTER/LAT_TIMR/T7 ;
  wire \MASTER/LAT_TIMR/T6 ;
  wire \MASTER/LAT_TIMR/OR_CE_L ;
  wire \MASTER/LAT_TIMR/T5 ;
  wire \MASTER/LAT_TIMR/T4 ;
  wire \MASTER/LAT_TIMR/$1I129/$1N2216 ;
  wire \MASTER/LAT_TIMR/Q4/TQ ;
  wire \MASTER/LAT_TIMR/Q4/MD ;
  wire \MASTER/LAT_TIMR/Q4/$1I30/M1 ;
  wire \MASTER/LAT_TIMR/Q4/$1I30/M0 ;
  wire \MASTER/LAT_TIMR/Q6/TQ ;
  wire \MASTER/LAT_TIMR/Q6/MD ;
  wire \MASTER/LAT_TIMR/Q6/$1I30/M1 ;
  wire \MASTER/LAT_TIMR/Q6/$1I30/M0 ;
  wire \MASTER/LAT_TIMR/Q7/TQ ;
  wire \MASTER/LAT_TIMR/Q7/MD ;
  wire \MASTER/LAT_TIMR/Q7/$1I30/M1 ;
  wire \MASTER/LAT_TIMR/Q7/$1I30/M0 ;
  wire \MASTER/LAT_TIMR/TIME_OUT/$1N2215 ;
  wire \MASTER/LAT_TIMR/TIME_OUT/D ;
  wire \MASTER/LAT_TIMR/Q5/TQ ;
  wire \MASTER/LAT_TIMR/Q5/MD ;
  wire \MASTER/LAT_TIMR/Q5/$1I30/M1 ;
  wire \MASTER/LAT_TIMR/Q5/$1I30/M0 ;
  wire \MASTER/LAT_TIMR/$2I121/$1N2216 ;
  wire \MASTER/LAT_TIMR/Q1/TQ ;
  wire \MASTER/LAT_TIMR/Q1/MD ;
  wire \MASTER/LAT_TIMR/Q1/$1I30/M1 ;
  wire \MASTER/LAT_TIMR/Q1/$1I30/M0 ;
  wire \MASTER/LAT_TIMR/Q0/TQ ;
  wire \MASTER/LAT_TIMR/Q0/MD ;
  wire \MASTER/LAT_TIMR/Q0/$1I30/M1 ;
  wire \MASTER/LAT_TIMR/Q0/$1I30/M0 ;
  wire \MASTER/LAT_TIMR/Q2/TQ ;
  wire \MASTER/LAT_TIMR/Q2/MD ;
  wire \MASTER/LAT_TIMR/Q2/$1I30/M1 ;
  wire \MASTER/LAT_TIMR/Q2/$1I30/M0 ;
  wire \MASTER/LAT_TIMR/Q3/TQ ;
  wire \MASTER/LAT_TIMR/Q3/MD ;
  wire \MASTER/LAT_TIMR/Q3/$1I30/M1 ;
  wire \MASTER/LAT_TIMR/Q3/$1I30/M0 ;
  wire \MASTER/PCI-0CH/$1N2518 ;
  wire \MASTER/PCI-0CH/$1N2513 ;
  wire \MASTER/$4I3254/$1N2216 ;
  wire \MASTER/$4I3319/$1N2216 ;
  wire \PCI-CNTL/NS_PWIN64 ;
  wire \PCI-CNTL/ANY_NS_BH64 ;
  wire \PCI-CNTL/ANY_BH64 ;
  wire \PCI-CNTL/$4N752 ;
  wire \PCI-CNTL/NS_CYC64 ;
  wire \PCI-CNTL/HOLDCYC ;
  wire \PCI-CNTL/NS_PWIN ;
  wire \PCI-CNTL/WIN_3628 ;
  wire \PCI-CNTL/TACK64- ;
  wire \PCI-CNTL/TSTOP- ;
  wire \PCI-CNTL/$1N1000 ;
  wire \PCI-CNTL/$1N988 ;
  wire \PCI-CNTL/TTRDY- ;
  wire \PCI-CNTL/TDEVSEL- ;
  wire \PCI-CNTL/CBE_N3 ;
  wire \PCI-CNTL/CBE_N2 ;
  wire \PCI-CNTL/CBE_N1 ;
  wire \PCI-CNTL/CBE_N0 ;
  wire \PCI-CNTL/DSTR ;
  wire \PCI-CNTL/END ;
  wire \PCI-CNTL/CMD15 ;
  wire \PCI-CNTL/CMD14 ;
  wire \PCI-CNTL/CMD13 ;
  wire \PCI-CNTL/CMD12 ;
  wire \PCI-CNTL/CMD11 ;
  wire \PCI-CNTL/CMD10 ;
  wire \PCI-CNTL/CMD9 ;
  wire \PCI-CNTL/CMD8 ;
  wire \PCI-CNTL/CMD7 ;
  wire \PCI-CNTL/CMD6 ;
  wire \PCI-CNTL/CMD5 ;
  wire \PCI-CNTL/CMD4 ;
  wire \PCI-CNTL/CMD3 ;
  wire \PCI-CNTL/CMD2 ;
  wire \PCI-CNTL/CMD1 ;
  wire \PCI-CNTL/CMD0 ;
  wire \PCI-CNTL/NS_CFG_HIT ;
  wire \PCI-CNTL/CFG_CYC ;
  wire \PCI-CNTL/LADX9 ;
  wire \PCI-CNTL/LADX8 ;
  wire \PCI-CNTL/LADX7 ;
  wire \PCI-CNTL/LADX6 ;
  wire \PCI-CNTL/LADX5 ;
  wire \PCI-CNTL/LADX4 ;
  wire \PCI-CNTL/LADX3 ;
  wire \PCI-CNTL/ADX15 ;
  wire \PCI-CNTL/LADX2 ;
  wire \PCI-CNTL/ADX14 ;
  wire \PCI-CNTL/LADX1 ;
  wire \PCI-CNTL/ADX13 ;
  wire \PCI-CNTL/LADX0 ;
  wire \PCI-CNTL/ADX12 ;
  wire \PCI-CNTL/ADX11 ;
  wire \PCI-CNTL/ADX10 ;
  wire \PCI-CNTL/LADX15 ;
  wire \PCI-CNTL/LADX14 ;
  wire \PCI-CNTL/LADX13 ;
  wire \PCI-CNTL/LADX12 ;
  wire \PCI-CNTL/LADX11 ;
  wire \PCI-CNTL/LADX10 ;
  wire \PCI-CNTL/ADX9 ;
  wire \PCI-CNTL/ADX8 ;
  wire \PCI-CNTL/ADX7 ;
  wire \PCI-CNTL/ADX6 ;
  wire \PCI-CNTL/ADX5 ;
  wire \PCI-CNTL/ADX4 ;
  wire \PCI-CNTL/ADX3 ;
  wire \PCI-CNTL/ADX2 ;
  wire \PCI-CNTL/ADX1 ;
  wire \PCI-CNTL/ADX0 ;
  wire \PCI-CNTL/S_ABORT ;
  wire \PCI-CNTL/HOLD_APERR ;
  wire \PCI-CNTL/PCI-LA/AD7610-0000 ;
  wire \PCI-CNTL/PCI-LA/$1N2762 ;
  wire \PCI-CNTL/PCI-LA/$1N2666 ;
  wire \PCI-CNTL/PCI-LA/$1N2668 ;
  wire \PCI-CNTL/PCI-LA/$1N2764 ;
  wire \PCI-CNTL/PCI-LA/$1N2670 ;
  wire \PCI-CNTL/PCI-LA/$1N2766 ;
  wire \PCI-CNTL/PCI-LA/$1N2672 ;
  wire \PCI-CNTL/PCI-LA/$1N2768 ;
  wire \PCI-CNTL/PCI-LA/$1N2760 ;
  wire \PCI-CNTL/PCI-LA/$1N2625 ;
  wire \PCI-CNTL/PCI-LA/$1N2620 ;
  wire \PCI-CNTL/PCI-LA/$1N2621 ;
  wire \PCI-CNTL/PCI-LA/$1N2619 ;
  wire \PCI-CNTL/PCI-LA/$1N2756 ;
  wire \PCI-CNTL/PCI-LA/$1N2623 ;
  wire \PCI-CNTL/PCI-LA/$1N2624 ;
  wire \PCI-CNTL/PCI-LA/DEC-A/$1N2277 ;
  wire \PCI-CNTL/PCI-LA/DEC-A/$1N2275 ;
  wire \PCI-CNTL/PCI-LA/DEC-B/$1N2277 ;
  wire \PCI-CNTL/PCI-LA/DEC-C/$1N2290 ;
  wire \PCI-CNTL/PCI-LA/DEC-C/$1N2289 ;
  wire \PCI-CNTL/PCI-LA/DEC-D/$1N2290 ;
  wire \PCI-CNTL/PCI-LA/DEC-E/$1N2275 ;
  wire \PCI-CNTL/PCI-LA/DEC-9/$1N2277 ;
  wire \PCI-CNTL/PCI-LA/DEC-9/$1N2276 ;
  wire \PCI-CNTL/PCI-LA/DEC-8/$1N2277 ;
  wire \PCI-CNTL/PCI-LA/DEC-8/$1N2276 ;
  wire \PCI-CNTL/PCI-LA/DEC-8/$1N2275 ;
  wire \PCI-CNTL/PCI-LA/DEC-7/$1N2283 ;
  wire \PCI-CNTL/PCI-LA/DEC-6/$1N2283 ;
  wire \PCI-CNTL/PCI-LA/DEC-6/$1N2275 ;
  wire \PCI-CNTL/PCI-LA/DEC-5/$1N2283 ;
  wire \PCI-CNTL/PCI-LA/DEC-5/$1N2276 ;
  wire \PCI-CNTL/PCI-LA/DEC-4/$1N2283 ;
  wire \PCI-CNTL/PCI-LA/DEC-4/$1N2276 ;
  wire \PCI-CNTL/PCI-LA/DEC-4/$1N2275 ;
  wire \PCI-CNTL/PCI-LA/DEC-3/$1N2283 ;
  wire \PCI-CNTL/PCI-LA/DEC-3/$1N2277 ;
  wire \PCI-CNTL/PCI-LA/DEC-2/$1N2283 ;
  wire \PCI-CNTL/PCI-LA/DEC-2/$1N2277 ;
  wire \PCI-CNTL/PCI-LA/DEC-2/$1N2275 ;
  wire \PCI-CNTL/PCI-LA/DEC-0/$1N2283 ;
  wire \PCI-CNTL/PCI-LA/DEC-0/$1N2277 ;
  wire \PCI-CNTL/PCI-LA/DEC-0/$1N2276 ;
  wire \PCI-CNTL/PCI-LA/DEC-0/$1N2275 ;
  wire \PCI-CNTL/PCI-LA/DEC-1/$1N2277 ;
  wire \PCI-CNTL/PCI-LA/DEC-1/$1N2278 ;
  wire \PCI-CNTL/PCI-LA/DEC-1/$1N2280 ;
  wire \PCI-CNTL/PCI-LA/0000/$1N2283 ;
  wire \PCI-CNTL/PCI-LA/0000/$1N2277 ;
  wire \PCI-CNTL/PCI-LA/0000/$1N2276 ;
  wire \PCI-CNTL/PCI-LA/0000/$1N2275 ;
  wire \PCI-CNTL/PCI-LC/$2N3210 ;
  wire \PCI-CNTL/PCI-LC/$2N3209 ;
  wire \PCI-CNTL/PCI-LC/TYPE00 ;
  wire \PCI-CNTL/PCI-LC/RW_CFG ;
  wire \PCI-CNTL/PCI-LC/NS_CFG_CYC ;
  wire \PCI-CNTL/PCI-LC/$2N2912 ;
  wire \PCI-CNTL/PCI-LC/DEC-E/$1N2275 ;
  wire \PCI-CNTL/PCI-LC/DEC-D/$1N2290 ;
  wire \PCI-CNTL/PCI-LC/DEC-C/$1N2290 ;
  wire \PCI-CNTL/PCI-LC/DEC-C/$1N2289 ;
  wire \PCI-CNTL/PCI-LC/DEC-0/$1N2283 ;
  wire \PCI-CNTL/PCI-LC/DEC-0/$1N2277 ;
  wire \PCI-CNTL/PCI-LC/DEC-0/$1N2276 ;
  wire \PCI-CNTL/PCI-LC/DEC-0/$1N2275 ;
  wire \PCI-CNTL/PCI-LC/DEC-1/$1N2277 ;
  wire \PCI-CNTL/PCI-LC/DEC-1/$1N2278 ;
  wire \PCI-CNTL/PCI-LC/DEC-1/$1N2280 ;
  wire \PCI-CNTL/PCI-LC/DEC-2/$1N2283 ;
  wire \PCI-CNTL/PCI-LC/DEC-2/$1N2277 ;
  wire \PCI-CNTL/PCI-LC/DEC-2/$1N2275 ;
  wire \PCI-CNTL/PCI-LC/DEC-3/$1N2283 ;
  wire \PCI-CNTL/PCI-LC/DEC-3/$1N2277 ;
  wire \PCI-CNTL/PCI-LC/DEC-4/$1N2283 ;
  wire \PCI-CNTL/PCI-LC/DEC-4/$1N2276 ;
  wire \PCI-CNTL/PCI-LC/DEC-4/$1N2275 ;
  wire \PCI-CNTL/PCI-LC/DEC-5/$1N2283 ;
  wire \PCI-CNTL/PCI-LC/DEC-5/$1N2276 ;
  wire \PCI-CNTL/PCI-LC/DEC-6/$1N2283 ;
  wire \PCI-CNTL/PCI-LC/DEC-6/$1N2275 ;
  wire \PCI-CNTL/PCI-LC/DEC-7/$1N2283 ;
  wire \PCI-CNTL/PCI-LC/DEC-8/$1N2277 ;
  wire \PCI-CNTL/PCI-LC/DEC-8/$1N2276 ;
  wire \PCI-CNTL/PCI-LC/DEC-8/$1N2275 ;
  wire \PCI-CNTL/PCI-LC/DEC-9/$1N2277 ;
  wire \PCI-CNTL/PCI-LC/DEC-9/$1N2276 ;
  wire \PCI-CNTL/PCI-LC/DEC-A/$1N2277 ;
  wire \PCI-CNTL/PCI-LC/DEC-A/$1N2275 ;
  wire \PCI-CNTL/PCI-LC/DEC-B/$1N2277 ;
  wire \PCI-CNTL/PCI-OE/UCS ;
  wire \PCI-CNTL/PCI-OE/$2N791 ;
  wire \PCI-CNTL/PCI-OE/LCS ;
  wire \PCI-CNTL/PCI-OE/$2N942 ;
  wire \PCI-CNTL/PCI-OE/00H ;
  wire \PCI-CNTL/PCI-OE/04H ;
  wire \PCI-CNTL/PCI-OE/08H ;
  wire \PCI-CNTL/PCI-OE/10H ;
  wire \PCI-CNTL/PCI-OE/14H ;
  wire \PCI-CNTL/PCI-OE/$2N744 ;
  wire \PCI-CNTL/PCI-OE/$2N745 ;
  wire \PCI-CNTL/PCI-OE/$2N746 ;
  wire \PCI-CNTL/PCI-OE/$2N747 ;
  wire \PCI-CNTL/PCI-OE/$2N748 ;
  wire \PCI-CNTL/PCI-OE/$2N749 ;
  wire \PCI-CNTL/PCI-OE/X ;
  wire \PCI-CNTL/PCI-OE/$2N750 ;
  wire \PCI-CNTL/PCI-OE/$2N751 ;
  wire \PCI-CNTL/PCI-OE/$2N752 ;
  wire \PCI-CNTL/PCI-OE/$2N753 ;
  wire \PCI-CNTL/PCI-OE/$2N754 ;
  wire \PCI-CNTL/PCI-OE/$2N755 ;
  wire \PCI-CNTL/PCI-OE/$2N756 ;
  wire \PCI-CNTL/PCI-OE/$2N757 ;
  wire \PCI-CNTL/PCI-OE/$2N758 ;
  wire \PCI-CNTL/PCI-OE/$2N697 ;
  wire \PCI-CNTL/PCI-OE/NS_OE_ROM ;
  wire \PCI-CNTL/PCI-OE/$2N795 ;
  wire \PCI-CNTL/PCI-OE/0CH ;
  wire \PCI-CNTL/PCI-OE/28H ;
  wire \PCI-CNTL/PCI-OE/2CH ;
  wire \PCI-CNTL/PCI-OE/18H ;
  wire \PCI-CNTL/PCI-OE/1CH ;
  wire \PCI-CNTL/PCI-OE/20H ;
  wire \PCI-CNTL/PCI-OE/24H ;
  wire \PCI-CNTL/PCI-OE/30H ;
  wire \PCI-CNTL/PCI-OE/34H ;
  wire \PCI-CNTL/PCI-OE/38H ;
  wire \PCI-CNTL/PCI-OE/3CH ;
  wire \PCI-CNTL/PCI-OE/OE15/R ;
  wire \PCI-CNTL/PCI-OE/OE15/$1N301 ;
  wire \PCI-CNTL/PCI-OE/OE15/S ;
  wire \PCI-CNTL/PCI-OE/OE15/Q ;
  wire \PCI-CNTL/PCI-OE/OE15/D ;
  wire \PCI-CNTL/PCI-OE/OE15/C ;
  wire \PCI-CNTL/PCI-OE/OE15/NS_OE ;
  wire \PCI-CNTL/PCI-OE/OE7/R ;
  wire \PCI-CNTL/PCI-OE/OE7/$1N301 ;
  wire \PCI-CNTL/PCI-OE/OE7/S ;
  wire \PCI-CNTL/PCI-OE/OE7/Q ;
  wire \PCI-CNTL/PCI-OE/OE7/D ;
  wire \PCI-CNTL/PCI-OE/OE7/C ;
  wire \PCI-CNTL/PCI-OE/OE7/NS_OE ;
  wire \PCI-CNTL/PCI-OE/OE6/R ;
  wire \PCI-CNTL/PCI-OE/OE6/$1N301 ;
  wire \PCI-CNTL/PCI-OE/OE6/S ;
  wire \PCI-CNTL/PCI-OE/OE6/Q ;
  wire \PCI-CNTL/PCI-OE/OE6/D ;
  wire \PCI-CNTL/PCI-OE/OE6/C ;
  wire \PCI-CNTL/PCI-OE/OE6/NS_OE ;
  wire \PCI-CNTL/PCI-OE/OE5/R ;
  wire \PCI-CNTL/PCI-OE/OE5/$1N301 ;
  wire \PCI-CNTL/PCI-OE/OE5/S ;
  wire \PCI-CNTL/PCI-OE/OE5/Q ;
  wire \PCI-CNTL/PCI-OE/OE5/D ;
  wire \PCI-CNTL/PCI-OE/OE5/C ;
  wire \PCI-CNTL/PCI-OE/OE5/NS_OE ;
  wire \PCI-CNTL/PCI-OE/OE4/R ;
  wire \PCI-CNTL/PCI-OE/OE4/$1N301 ;
  wire \PCI-CNTL/PCI-OE/OE4/S ;
  wire \PCI-CNTL/PCI-OE/OE4/Q ;
  wire \PCI-CNTL/PCI-OE/OE4/D ;
  wire \PCI-CNTL/PCI-OE/OE4/C ;
  wire \PCI-CNTL/PCI-OE/OE4/NS_OE ;
  wire \PCI-CNTL/PCI-OE/OE3/R ;
  wire \PCI-CNTL/PCI-OE/OE3/$1N301 ;
  wire \PCI-CNTL/PCI-OE/OE3/S ;
  wire \PCI-CNTL/PCI-OE/OE3/Q ;
  wire \PCI-CNTL/PCI-OE/OE3/D ;
  wire \PCI-CNTL/PCI-OE/OE3/C ;
  wire \PCI-CNTL/PCI-OE/OE3/NS_OE ;
  wire \PCI-CNTL/PCI-OE/OE8/R ;
  wire \PCI-CNTL/PCI-OE/OE8/$1N301 ;
  wire \PCI-CNTL/PCI-OE/OE8/S ;
  wire \PCI-CNTL/PCI-OE/OE8/Q ;
  wire \PCI-CNTL/PCI-OE/OE8/D ;
  wire \PCI-CNTL/PCI-OE/OE8/C ;
  wire \PCI-CNTL/PCI-OE/OE8/NS_OE ;
  wire \PCI-CNTL/PCI-OE/OE9/R ;
  wire \PCI-CNTL/PCI-OE/OE9/$1N301 ;
  wire \PCI-CNTL/PCI-OE/OE9/S ;
  wire \PCI-CNTL/PCI-OE/OE9/Q ;
  wire \PCI-CNTL/PCI-OE/OE9/D ;
  wire \PCI-CNTL/PCI-OE/OE9/C ;
  wire \PCI-CNTL/PCI-OE/OE9/NS_OE ;
  wire \PCI-CNTL/PCI-OE/OE12/R ;
  wire \PCI-CNTL/PCI-OE/OE12/$1N301 ;
  wire \PCI-CNTL/PCI-OE/OE12/S ;
  wire \PCI-CNTL/PCI-OE/OE12/Q ;
  wire \PCI-CNTL/PCI-OE/OE12/D ;
  wire \PCI-CNTL/PCI-OE/OE12/C ;
  wire \PCI-CNTL/PCI-OE/OE12/NS_OE ;
  wire \PCI-CNTL/PCI-OE/OE1/R ;
  wire \PCI-CNTL/PCI-OE/OE1/$1N301 ;
  wire \PCI-CNTL/PCI-OE/OE1/S ;
  wire \PCI-CNTL/PCI-OE/OE1/Q ;
  wire \PCI-CNTL/PCI-OE/OE1/D ;
  wire \PCI-CNTL/PCI-OE/OE1/C ;
  wire \PCI-CNTL/PCI-OE/OE1/NS_OE ;
  wire \PCI-CNTL/PCI-OE/$1I849/$1N2216 ;
  wire \PCI-CNTL/PCI-OE/$1I850/$1N2216 ;
  wire \PCI-CNTL/PCI-OE/$1I853/$1N2216 ;
  wire \PCI-CNTL/PCI-OE/$1I868/$1N2216 ;
  wire \PCI-CNTL/PCI-OE/$1I870/$1N2216 ;
  wire \PCI-CNTL/PCI-OE/$1I872/$1N2216 ;
  wire \PCI-CNTL/PCI-OE/DEC-E/$1N2275 ;
  wire \PCI-CNTL/PCI-OE/DEC-D/$1N2290 ;
  wire \PCI-CNTL/PCI-OE/DEC-C/$1N2290 ;
  wire \PCI-CNTL/PCI-OE/DEC-C/$1N2289 ;
  wire \PCI-CNTL/PCI-OE/DEC-9/$1N2277 ;
  wire \PCI-CNTL/PCI-OE/DEC-9/$1N2276 ;
  wire \PCI-CNTL/PCI-OE/DEC-8/$1N2277 ;
  wire \PCI-CNTL/PCI-OE/DEC-8/$1N2276 ;
  wire \PCI-CNTL/PCI-OE/DEC-8/$1N2275 ;
  wire \PCI-CNTL/PCI-OE/DEC-7/$1N2283 ;
  wire \PCI-CNTL/PCI-OE/DEC-6/$1N2283 ;
  wire \PCI-CNTL/PCI-OE/DEC-6/$1N2275 ;
  wire \PCI-CNTL/PCI-OE/DEC-B/$1N2277 ;
  wire \PCI-CNTL/PCI-OE/DEC-A/$1N2277 ;
  wire \PCI-CNTL/PCI-OE/DEC-A/$1N2275 ;
  wire \PCI-CNTL/PCI-OE/DEC-3/$1N2283 ;
  wire \PCI-CNTL/PCI-OE/DEC-3/$1N2277 ;
  wire \PCI-CNTL/PCI-OE/$2I617/D ;
  wire \PCI-CNTL/PCI-OE/$2I617/$1N18 ;
  wire \PCI-CNTL/PCI-OE/OR16/$1N2234 ;
  wire \PCI-CNTL/PCI-OE/OR16/$1N2243 ;
  wire \PCI-CNTL/PCI-OE/OR16/$1N2224 ;
  wire \PCI-CNTL/PCI-OE/OR16/$1N2216 ;
  wire \PCI-CNTL/PCI-OE/DEC-5/$1N2283 ;
  wire \PCI-CNTL/PCI-OE/DEC-5/$1N2276 ;
  wire \PCI-CNTL/PCI-OE/DEC-4/$1N2283 ;
  wire \PCI-CNTL/PCI-OE/DEC-4/$1N2276 ;
  wire \PCI-CNTL/PCI-OE/DEC-4/$1N2275 ;
  wire \PCI-CNTL/PCI-OE/DEC-2/$1N2283 ;
  wire \PCI-CNTL/PCI-OE/DEC-2/$1N2277 ;
  wire \PCI-CNTL/PCI-OE/DEC-2/$1N2275 ;
  wire \PCI-CNTL/PCI-OE/DEC-1/$1N2277 ;
  wire \PCI-CNTL/PCI-OE/DEC-1/$1N2278 ;
  wire \PCI-CNTL/PCI-OE/DEC-1/$1N2280 ;
  wire \PCI-CNTL/PCI-OE/DEC-0/$1N2283 ;
  wire \PCI-CNTL/PCI-OE/DEC-0/$1N2277 ;
  wire \PCI-CNTL/PCI-OE/DEC-0/$1N2276 ;
  wire \PCI-CNTL/PCI-OE/DEC-0/$1N2275 ;
  wire \PCI-CNTL/PCI-OE/SW1/$1I2290/$1N2216 ;
  wire \PCI-CNTL/PCI-OE/SW15/$1I2290/$1N2216 ;
  wire \PCI-CNTL/PCI-OE/SW3/$1I2290/$1N2216 ;
  wire \PCI-CNTL/$1I995/$1N2215 ;
  wire \PCI-CNTL/$1I995/D ;
  wire \PCI-CNTL/PCI-TSM/PCI-IDLE/BKOF_NS_TNAR ;
  wire \PCI-CNTL/PCI-TSM/PCI-IDLE/DATA_NS_TNAR ;
  wire \PCI-CNTL/PCI-TSM/PCI-IDLE/EQN-A ;
  wire \PCI-CNTL/PCI-TSM/PCI-IDLE/$1N483 ;
  wire \PCI-CNTL/PCI-TSM/PCI-IDLE/$1N367 ;
  wire \PCI-CNTL/PCI-TSM/PCI-IDLE/NS_TNAR ;
  wire \PCI-CNTL/PCI-TSM/PCI-IDLE/IDLE_NS_IDLE ;
  wire \PCI-CNTL/PCI-TSM/PCI-IDLE/BUSY_NS_IDLE ;
  wire \PCI-CNTL/PCI-TSM/PCI-IDLE/NS_IDLE ;
  wire \PCI-CNTL/PCI-TSM/PCI-BUSY/BUSY_NS_BUSY ;
  wire \PCI-CNTL/PCI-TSM/PCI-BUSY/NS_BUSY ;
  wire \PCI-CNTL/PCI-TSM/PCI-BUSY/IDLE_NS_BUSY ;
  wire \PCI-CNTL/PCI-TSM/PCI-BUSY/HITIDLEORBUSY ;
  wire \PCI-CNTL/PCI-TSM/PCI-BUSY/$1N484 ;
  wire \PCI-CNTL/PCI-TSM/PCI-BUSY/$1N476 ;
  wire \PCI-CNTL/PCI-TSM/PCI-BUSY/EQN-B ;
  wire \PCI-CNTL/PCI-TSM/PCI-BUSY/EQN-A ;
  wire \PCI-CNTL/PCI-TSM/PCI-DATA/$1N673 ;
  wire \PCI-CNTL/PCI-TSM/PCI-DATA/EQN-B ;
  wire \PCI-CNTL/PCI-TSM/PCI-DATA/$1N628 ;
  wire \PCI-CNTL/PCI-TSM/PCI-DATA/CBUSY_NS_DATA ;
  wire \PCI-CNTL/PCI-TSM/PCI-DATA/NS_DATA ;
  wire \PCI-CNTL/PCI-TSM/PCI-DATA/DATA_NS_DATA ;
  wire \PCI-CNTL/PCI-TSM/PCI-DATA/EQN-E ;
  wire \PCI-CNTL/PCI-TSM/PCI-DATA/$1N497 ;
  wire \PCI-CNTL/PCI-TSM/PCI-DATA/$1N483 ;
  wire \PCI-CNTL/PCI-TSM/PCI-DATA/$1N495 ;
  wire \PCI-CNTL/PCI-TSM/PCI-DATA/BUSY_NS_DATA ;
  wire \PCI-CNTL/PCI-TSM/PCI-DATA/EQN-A ;
  wire \PCI-CNTL/PCI-TSM/PCI-DATA/HIT ;
  wire \PCI-CNTL/PCI-TSM/PCI-DATA/EQN-D ;
  wire \PCI-CNTL/PCI-TSM/PCI-DATA/$1N452 ;
  wire \PCI-CNTL/PCI-TSM/PCI-BKOF/EQN-AB ;
  wire \PCI-CNTL/PCI-TSM/PCI-BKOF/BKOF_HIT ;
  wire \PCI-CNTL/PCI-TSM/PCI-BKOF/S_EQN ;
  wire \PCI-CNTL/PCI-TSM/PCI-BKOF/C_EQN ;
  wire \PCI-CNTL/PCI-TSM/PCI-BKOF/EQN-B ;
  wire \PCI-CNTL/PCI-TSM/PCI-BKOF/$1N531 ;
  wire \PCI-CNTL/PCI-TSM/PCI-BKOF/IDLE_BUSY_NS ;
  wire \PCI-CNTL/PCI-TSM/PCI-BKOF/HIT ;
  wire \PCI-CNTL/PCI-TSM/PCI-BKOF/EQN-E ;
  wire \PCI-CNTL/PCI-TSM/PCI-BKOF/$1N479 ;
  wire \PCI-CNTL/PCI-TSM/PCI-BKOF/$1N477 ;
  wire \PCI-CNTL/PCI-TSM/PCI-BKOF/EQN-A ;
  wire \PCI-CNTL/PCI-TSM/PCI-BKOF/TURNIDLE ;
  wire \PCI-CNTL/PCI-TSM/PCI-BKOF/DATA_NS ;
  wire \PCI-CNTL/PCI-TSM/PCI-BKOF/DATA_NS_BKOF ;
  wire \PCI-CNTL/PCI-TSM/PCI-BKOF/BKOF_NS_BKOF ;
  wire \PCI-CNTL/PCI-TSM/PCI-BKOF/NS_BKOF ;
  wire \PCI-CNTL/PCI-TSM/$1I426/$1N2216 ;
  wire \PCI-CNTL/PCI-OFCN/HIT ;
  wire \PCI-CNTL/PCI-OFCN/NL_MEM ;
  wire \PCI-CNTL/PCI-OFCN/$1N1433 ;
  wire \PCI-CNTL/PCI-OFCN/$1N1431 ;
  wire \PCI-CNTL/PCI-OFCN/ACKHIT ;
  wire \PCI-CNTL/PCI-OFCN/PCI-AK64/$3N836 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-AK64/NS_F0 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-AK64/$2N969 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-AK64/$2N970 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-AK64/$2N974 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-AK64/$2N968 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-AK64/$2N982 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-AK64/$2N962 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-AK64/$2N931 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-AK64/$2N937 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-AK64/NS_F0_I1 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-AK64/DUCKLING ;
  wire \PCI-CNTL/PCI-OFCN/PCI-AK64/NS_F0_I0 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-AK64/DATA_NS_DATA_OR_BKOF0 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-AK64/BKOF_NS_BKOF ;
  wire \PCI-CNTL/PCI-OFCN/PCI-AK64/DATA_NS_DATA_OR_BKOF1 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-AK64/EQN-F1A ;
  wire \PCI-CNTL/PCI-OFCN/PCI-AK64/EQN-C ;
  wire \PCI-CNTL/PCI-OFCN/PCI-AK64/NS_HIT ;
  wire \PCI-CNTL/PCI-OFCN/PCI-AK64/$1N809 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-AK64/$1N794 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-AK64/$1N795 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-AK64/$1N789 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-AK64/NS_F1 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-AK64/LATE_GATE ;
  wire \PCI-CNTL/PCI-OFCN/PCI-AK64/$1N801 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-AK64/$1N846 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-AK64/$1N782 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-AK64/$3I854/M1 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-AK64/$3I854/M0 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-AK64/$3I864/$1N2216 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-DSEL/$3N806 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-DSEL/NS_F0 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-DSEL/$2N972 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-DSEL/$2N979 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-DSEL/$2N938 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-DSEL/$2N939 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-DSEL/$2N899 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-DSEL/NS_F0_I0 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-DSEL/$2N917 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-DSEL/NS_F0_I1 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-DSEL/DATA_NS_DATA_OR_BKOF1 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-DSEL/BKOF_NS_BKOF ;
  wire \PCI-CNTL/PCI-OFCN/PCI-DSEL/$2N875 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-DSEL/$2N893 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-DSEL/DUCKLING ;
  wire \PCI-CNTL/PCI-OFCN/PCI-DSEL/DATA_NS_DATA_OR_BKOF0 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-DSEL/$1N784 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-DSEL/$1N923 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-DSEL/$1N783 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-DSEL/$1N790 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-DSEL/NS_F1 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-DSEL/LATE_GATE ;
  wire \PCI-CNTL/PCI-OFCN/PCI-DSEL/$1N919 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-DSEL/EQN-F1A ;
  wire \PCI-CNTL/PCI-OFCN/PCI-DSEL/EQN-C ;
  wire \PCI-CNTL/PCI-OFCN/PCI-DSEL/$1N1033 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-DSEL/$1N1030 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-DSEL/NS_HIT ;
  wire \PCI-CNTL/PCI-OFCN/PCI-DSEL/$3I798/M1 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-DSEL/$3I798/M0 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-DSEL/$3I813/$1N2216 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-TRDY/S_FIRSTIN ;
  wire \PCI-CNTL/PCI-OFCN/PCI-TRDY/$4N968 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-TRDY/$4N1042 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-TRDY/$4N1052 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-TRDY/S_FIRST0 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-TRDY/SF0_I1 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-TRDY/SF0_I0 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-TRDY/$4N1030 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-TRDY/$4N1002 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-TRDY/S_FIRST1 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-TRDY/$4N1008 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-TRDY/TRDY_OFF ;
  wire \PCI-CNTL/PCI-OFCN/PCI-TRDY/$3N833 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-TRDY/$3N837 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-TRDY/$3N835 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-TRDY/HOLD_TRDY ;
  wire \PCI-CNTL/PCI-OFCN/PCI-TRDY/SWAN1 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-TRDY/SWAN2 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-TRDY/$1N786 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-TRDY/SWAN0 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-TRDY/$1N763 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-TRDY/NS_TRDY- ;
  wire \PCI-CNTL/PCI-OFCN/PCI-TRDY/CRABILL ;
  wire \PCI-CNTL/PCI-OFCN/PCI-TRDY/BUSY_NS_DATA ;
  wire \PCI-CNTL/PCI-OFCN/PCI-TRDY/C_EQN ;
  wire \PCI-CNTL/PCI-OFCN/PCI-TRDY/$1N738 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-TRDY/$1N735 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-TRDY/S_EQN ;
  wire \PCI-CNTL/PCI-OFCN/PCI-TRDY/HIT ;
  wire \PCI-CNTL/PCI-OFCN/PCI-TRDY/EQN-A ;
  wire \PCI-CNTL/PCI-OFCN/PCI-TRDY/DATA_NS_DATA ;
  wire \PCI-CNTL/PCI-OFCN/PCI-TRDY/EQN-F ;
  wire \PCI-CNTL/PCI-OFCN/PCI-TRDY/EQN-E ;
  wire \PCI-CNTL/PCI-OFCN/PCI-TRDY/$1N497 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-TRDY/$1N637 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-TRDY/$1N495 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-TRDY/$1N466 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-TRDY/EQN-D ;
  wire \PCI-CNTL/PCI-OFCN/PCI-TRDY/$1N452 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I782/M1 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I782/M0 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-TRDY/$3I957/$1N2216 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-TRDY/$4I1028/M1 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-TRDY/$4I1028/M0 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-STOP/NS_1 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-STOP/$3N1288 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-STOP/$3N1280 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-STOP/$3N1277 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-STOP/NS_0 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-STOP/$3N1256 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-STOP/$3N1259 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-STOP/$3N1257 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-STOP/$1N1503 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-STOP/$1N1500 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-STOP/SUB_DATA ;
  wire \PCI-CNTL/PCI-OFCN/PCI-STOP/$1N1459 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-STOP/PRE_NS ;
  wire \PCI-CNTL/PCI-OFCN/PCI-STOP/$1N1453 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-STOP/$1N1434 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-STOP/$1N1438 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-STOP/I_DATA_FLAG ;
  wire \PCI-CNTL/PCI-OFCN/PCI-STOP/TERM_OTHER ;
  wire \PCI-CNTL/PCI-OFCN/PCI-STOP/TERM ;
  wire \PCI-CNTL/PCI-OFCN/PCI-STOP/DIS_WDATA ;
  wire \PCI-CNTL/PCI-OFCN/PCI-STOP/HIT ;
  wire \PCI-CNTL/PCI-OFCN/PCI-STOP/PRE_DATA ;
  wire \PCI-CNTL/PCI-OFCN/PCI-STOP/TERMINATE ;
  wire \PCI-CNTL/PCI-OFCN/PCI-STOP/$1N1266 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-STOP/IDATA_WIN ;
  wire \PCI-CNTL/PCI-OFCN/PCI-STOP/FAST_TERM_WIN ;
  wire \PCI-CNTL/PCI-OFCN/PCI-STOP/PRE_DEVSEL ;
  wire \PCI-CNTL/PCI-OFCN/PCI-STOP/$1N1159 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-STOP/JAYANT ;
  wire \PCI-CNTL/PCI-OFCN/PCI-STOP/NUPUR ;
  wire \PCI-CNTL/PCI-OFCN/PCI-STOP/WR_OR_NRDY ;
  wire \PCI-CNTL/PCI-OFCN/PCI-STOP/READY ;
  wire \PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1368/M1 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1368/M0 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1373/M1 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1373/M0 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1437/$1N2215 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1437/D ;
  wire \PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1499/M1 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1499/M0 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-STOP/$3I1332/$1N2216 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/SET_LB64 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/SET_LT64 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/SET_T64 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/SET_B64 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/NS-OE_ADO_B64 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/NS-OE_ADO_T64 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/NS-OE_ADO_LB64 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/NS-OE_ADO_LT64 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/EQN-D64 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/$5N1020 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/$5N1019 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/$5N1023 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/$5N1033 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/BH64_012 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/BEGIN64 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/B_BUSY_NS64 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/S_EQN64 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/END64 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/TRSTOPQ64 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/SET_LB ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/SET_LT ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/SET_T ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/SET_B ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/NS-OE_ADO_B ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/NS-OE_ADO_T ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/NS-OE_ADO_LB ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/NS-OE_ADO_LT ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/BEGIN ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/$3N905 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/$3N903 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/$3N918 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/C_EQN ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/B_BUSY_NS ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/$3N893 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/END ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/$3N861 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/TRSTOPQ ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/$3N818 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/S_EQN ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/BHIT_012 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/EQN-D ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/$3N628 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/$2N1335 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/ACTIVE64 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/NS_HIT64 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/$2N1272 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/OE_ACK64_IN ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/$2N1220 ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/NS_HIT ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/OE_TRDY_IN ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/ACTIVE ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/HOLD_OE_PERR ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/SET_OE_PERR ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/TRDYDEL ;
  wire \PCI-CNTL/PCI-OFCN/PCI-XOE/EQN-A ;
  wire \PCI-CNTL/$4I614/M1 ;
  wire \PCI-CNTL/$4I614/M0 ;
  wire \TDLY/$1N332 ;
  wire \TDLY/$1N318 ;
  wire \TDLY/D6_4118 ;
  wire \TDLY/D5_4117 ;
  wire \TDLY/D4_4116 ;
  wire \TDLY/D3_4115 ;
  wire \TDLY/D2_4114 ;
  wire \TDLY/D1_4113 ;
  wire \TDLY/$1I315/M23 ;
  wire \TDLY/$1I315/M01 ;
  wire \TDLY/$1I315/M01/M0 ;
  wire \TDLY/$1I315/M01/M1 ;
  wire \TDLY/$1I315/M23/M0 ;
  wire \TDLY/$1I315/M23/M1 ;
  wire \TDLY/$1I319/$1N2216 ;
  wire \TDLY/$1I328/M23 ;
  wire \TDLY/$1I328/M01 ;
  wire \TDLY/$1I328/M01/M0 ;
  wire \TDLY/$1I328/M01/M1 ;
  wire \TDLY/$1I328/M23/M0 ;
  wire \TDLY/$1I328/M23/M1 ;
  wire \TDLY/$1I331/$1N2216 ;
  wire \IDLY/$1N332 ;
  wire \IDLY/$1N318 ;
  wire \IDLY/D6_4183 ;
  wire \IDLY/D5_4182 ;
  wire \IDLY/D4_4181 ;
  wire \IDLY/D3_4180 ;
  wire \IDLY/D2_4179 ;
  wire \IDLY/D1_4178 ;
  wire \IDLY/$1I315/M23 ;
  wire \IDLY/$1I315/M01 ;
  wire \IDLY/$1I315/M01/M0 ;
  wire \IDLY/$1I315/M01/M1 ;
  wire \IDLY/$1I315/M23/M0 ;
  wire \IDLY/$1I315/M23/M1 ;
  wire \IDLY/$1I319/$1N2216 ;
  wire \IDLY/$1I328/M23 ;
  wire \IDLY/$1I328/M01 ;
  wire \IDLY/$1I328/M01/M0 ;
  wire \IDLY/$1I328/M01/M1 ;
  wire \IDLY/$1I328/M23/M0 ;
  wire \IDLY/$1I328/M23/M1 ;
  wire \IDLY/$1I331/$1N2216 ;
  wire \DATA_VLD/NS_SDV ;
  wire \DATA_VLD/NS_MDV ;
  wire \SRC_EN/MDATA_EQN ;
  wire \SRC_EN/S_SRC_PRE ;
  wire \SRC_EN/SFIRST_EQN ;
  wire \SRC_EN/SDATA_EQN ;
  wire \OUT_CE/HARD_CE ;
  wire \OUT_CE/$3N1089 ;
  wire \OUT_CE/$3N1090 ;
  wire \OUT_CE/FIRST ;
  wire \OUT_CE/$3N1041 ;
  wire \OUT_CE/SOFT_CE ;
  wire \OUT_CE/M_CE_XX0 ;
  wire \OUT_CE/M_CE_XX1 ;
  wire \OUT_CE/$2N1066 ;
  wire \OUT_CE/$2N1067 ;
  wire \OUT_CE/SOFT_CE0 ;
  wire \OUT_CE/S_CE_XX0 ;
  wire \OUT_CE/SOFT_CE1 ;
  wire \OUT_CE/S_CE_XX1 ;
  wire \OUT_CE/M_CE_P1 ;
  wire \OUT_CE/M_OK_N ;
  wire \OUT_CE/$2N1025 ;
  wire \OUT_CE/M_CE_P0 ;
  wire \OUT_CE/FFA_4285 ;
  wire \OUT_CE/S_CE_P0 ;
  wire \OUT_CE/NS_PAR_CE ;
  wire \OUT_CE/NS_PAR_CE1 ;
  wire \OUT_CE/NS_PAR_CE0 ;
  wire \OUT_CE/S_CE_P1 ;
  wire \OUT_CE/S_OK_N ;
  wire \OUT_CE/$2N1024 ;
  wire \OUT_CE/S_ND_T0 ;
  wire \OUT_CE/$1N989 ;
  wire \OUT_CE/MND_4275 ;
  wire \OUT_CE/$1N968 ;
  wire \OUT_CE/S_ND_T1 ;
  wire \OUT_CE/NS_NEWDATA ;
  wire \OUT_CE/ZERO_ND_T1 ;
  wire \OUT_CE/M_ND_T1 ;
  wire \OUT_CE/ZERO_ND_T0 ;
  wire \OUT_CE/M_ND_T0 ;
  wire \OUT_CE/SND_4267 ;
  wire \OUT_CE/FANF_4266 ;
  wire \OUT_CE/$1I987/$1N2216 ;
  wire \OUT_CE/$1I988/$1N2216 ;
  wire \OUT_CE/$2I1022/$1N2216 ;
  wire \OUT_CE/$2I1023/$1N2216 ;
  wire \OUT_CE/$2I1049/$1N2216 ;
  wire \OUT_CE/$2I1050/$1N2216 ;
  wire \OUT_CE/MAGICBOX/I3_NAND_TRDY_4239 ;
  wire \OUT_CE/MAGICBOX/I1_NAND_IRDY_4238 ;
  wire \OUT_CE/$4I1005/M1 ;
  wire \OUT_CE/$4I1005/M0 ;
  wire \OUT_SEL/$1N959 ;
  wire \OUT_SEL/$1N958 ;
  wire \OUT_SEL/SEL64_IN ;
  wire \OUT_SEL/$1N898 ;
  wire \OUT_SEL/$1N851 ;
  wire \OUT_SEL/S_IN ;
  wire \OUT_SEL/M_IN ;
  wire \OUT_SEL/$1N826 ;
  wire \OUT_SEL/$1N821 ;
  wire \OUT_SEL/$1N765 ;
  wire \OUT_SEL/$1N766 ;
  wire \OUT_SEL/SEL_IN ;
  wire \ADDR_VLD/$1N3964 ;
  wire \ADDR_VLD/TEMP_0 ;
  wire \ADDR_VLD/$1N3898 ;
  wire \ADDR_VLD/$1N3884 ;
  wire \ADDR_VLD/$1N3858 ;
  wire \ADDR_VLD/TEMP_1 ;
  wire \ADDR_VLD/TEMP_2 ;
  wire \ADDR_VLD/FRAMEQ- ;
  wire \ADDR_VLD/REQ64Q- ;
  wire \EOT/$1N630 ;
  wire \EOT/$1N631 ;
  wire \EOT/EQN-V1 ;
  wire \EOT/EQN-W1 ;
  wire \EOT/$1N627 ;
  wire \EOT/$1N623 ;
  wire \EOT/$1N624 ;
  wire \EOT/$1N658 ;
  wire \EOT/$1N603 ;
  wire \EOT/NS_1 ;
  wire \EOT/EOT_DL_4369 ;
  wire \EOT/EOT_D ;
  wire \EOT/NS_0 ;
  wire \EOT/EQN-W0 ;
  wire \EOT/EQN-V0 ;
  wire \PCI-PAR/PREP ;
  wire \PCI-PAR/$7N2995 ;
  wire \PCI-PAR/$7N2992 ;
  wire \PCI-PAR/PREN ;
  wire \PCI-PAR/PRE64N ;
  wire \PCI-PAR/PRE64P ;
  wire \PCI-PAR/X14O ;
  wire \PCI-PAR/DOQ59 ;
  wire \PCI-PAR/DOQ58 ;
  wire \PCI-PAR/DOQ57 ;
  wire \PCI-PAR/DOQ56 ;
  wire \PCI-PAR/X13O ;
  wire \PCI-PAR/DOQ55 ;
  wire \PCI-PAR/DOQ54 ;
  wire \PCI-PAR/DOQ53 ;
  wire \PCI-PAR/DOQ52 ;
  wire \PCI-PAR/X12O ;
  wire \PCI-PAR/DOQ51 ;
  wire \PCI-PAR/DOQ50 ;
  wire \PCI-PAR/DOQ49 ;
  wire \PCI-PAR/DOQ48 ;
  wire \PCI-PAR/X11O ;
  wire \PCI-PAR/DOQ47 ;
  wire \PCI-PAR/DOQ46 ;
  wire \PCI-PAR/DOQ45 ;
  wire \PCI-PAR/DOQ44 ;
  wire \PCI-PAR/X10O ;
  wire \PCI-PAR/DOQ43 ;
  wire \PCI-PAR/DOQ42 ;
  wire \PCI-PAR/DOQ41 ;
  wire \PCI-PAR/DOQ40 ;
  wire \PCI-PAR/X9O ;
  wire \PCI-PAR/DOQ39 ;
  wire \PCI-PAR/DOQ38 ;
  wire \PCI-PAR/DOQ37 ;
  wire \PCI-PAR/DOQ36 ;
  wire \PCI-PAR/X8O ;
  wire \PCI-PAR/DOQ35 ;
  wire \PCI-PAR/DOQ34 ;
  wire \PCI-PAR/DOQ33 ;
  wire \PCI-PAR/DOQ32 ;
  wire \PCI-PAR/X15O ;
  wire \PCI-PAR/DOQ63 ;
  wire \PCI-PAR/DOQ62 ;
  wire \PCI-PAR/DOQ61 ;
  wire \PCI-PAR/DOQ60 ;
  wire \PCI-PAR/AD_PAR64 ;
  wire \PCI-PAR/P7O ;
  wire \PCI-PAR/P6O ;
  wire \PCI-PAR/P5O ;
  wire \PCI-PAR/P4O ;
  wire \PCI-PAR/AD_PAR ;
  wire \PCI-PAR/P3O ;
  wire \PCI-PAR/P2O ;
  wire \PCI-PAR/P1O ;
  wire \PCI-PAR/P0O ;
  wire \PCI-PAR/X7O ;
  wire \PCI-PAR/DOQ31 ;
  wire \PCI-PAR/DOQ30 ;
  wire \PCI-PAR/DOQ29 ;
  wire \PCI-PAR/DOQ28 ;
  wire \PCI-PAR/X6O ;
  wire \PCI-PAR/DOQ27 ;
  wire \PCI-PAR/DOQ26 ;
  wire \PCI-PAR/DOQ25 ;
  wire \PCI-PAR/DOQ24 ;
  wire \PCI-PAR/X5O ;
  wire \PCI-PAR/DOQ23 ;
  wire \PCI-PAR/DOQ22 ;
  wire \PCI-PAR/DOQ21 ;
  wire \PCI-PAR/DOQ20 ;
  wire \PCI-PAR/X4O ;
  wire \PCI-PAR/DOQ19 ;
  wire \PCI-PAR/DOQ18 ;
  wire \PCI-PAR/DOQ17 ;
  wire \PCI-PAR/DOQ16 ;
  wire \PCI-PAR/X3O ;
  wire \PCI-PAR/DOQ15 ;
  wire \PCI-PAR/DOQ14 ;
  wire \PCI-PAR/DOQ13 ;
  wire \PCI-PAR/DOQ12 ;
  wire \PCI-PAR/X2O ;
  wire \PCI-PAR/DOQ11 ;
  wire \PCI-PAR/DOQ10 ;
  wire \PCI-PAR/DOQ9 ;
  wire \PCI-PAR/DOQ8 ;
  wire \PCI-PAR/X1O ;
  wire \PCI-PAR/DOQ7 ;
  wire \PCI-PAR/DOQ6 ;
  wire \PCI-PAR/DOQ5 ;
  wire \PCI-PAR/DOQ4 ;
  wire \PCI-PAR/X0O ;
  wire \PCI-PAR/DOQ3 ;
  wire \PCI-PAR/DOQ2 ;
  wire \PCI-PAR/DOQ1 ;
  wire \PCI-PAR/DOQ0 ;
  wire \PCI-PAR/PRE_APERR_N ;
  wire \PCI-PAR/$4N3107 ;
  wire \PCI-PAR/$4N3125 ;
  wire \PCI-PAR/PAP_0 ;
  wire \PCI-PAR/PAP32_0 ;
  wire \PCI-PAR/PAP64_0 ;
  wire \PCI-PAR/$4N3113 ;
  wire \PCI-PAR/CHECK64 ;
  wire \PCI-PAR/$4N3110 ;
  wire \PCI-PAR/CHECK32 ;
  wire \PCI-PAR/PAP_1 ;
  wire \PCI-PAR/PAP32_1 ;
  wire \PCI-PAR/PAP64_1 ;
  wire \PCI-PAR/$4N3109 ;
  wire \PCI-PAR/$4N3098 ;
  wire \PCI-PAR/M_DATAQ ;
  wire \PCI-PAR/$3N3054 ;
  wire \PCI-PAR/NS_1 ;
  wire \PCI-PAR/ERR32_1 ;
  wire \PCI-PAR/ERR64_1 ;
  wire \PCI-PAR/$3N3025 ;
  wire \PCI-PAR/$3N3024 ;
  wire \PCI-PAR/$3N3020 ;
  wire \PCI-PAR/NS_0 ;
  wire \PCI-PAR/$3N2935 ;
  wire \PCI-PAR/NS_SERR ;
  wire \PCI-PAR/$3N2930 ;
  wire \PCI-PAR/ADDR_VLDQ ;
  wire \PCI-PAR/NS_OE_SERR ;
  wire \PCI-PAR/ERR64_0 ;
  wire \PCI-PAR/PWIN64 ;
  wire \PCI-PAR/$3N2766 ;
  wire \PCI-PAR/ERR32_0 ;
  wire \PCI-PAR/PWIN ;
  wire \PCI-PAR/LC_PERR- ;
  wire \PCI-PAR/$3N2500 ;
  wire \PCI-PAR/$3N2761 ;
  wire \PCI-PAR/PER64_4858 ;
  wire \PCI-PAR/P7I ;
  wire \PCI-PAR/X15I ;
  wire \PCI-PAR/P6I ;
  wire \PCI-PAR/P5I ;
  wire \PCI-PAR/P4I ;
  wire \PCI-PAR/X8I ;
  wire \PCI-PAR/X9I ;
  wire \PCI-PAR/X11I ;
  wire \PCI-PAR/X10I ;
  wire \PCI-PAR/X12I ;
  wire \PCI-PAR/X13I ;
  wire \PCI-PAR/X14I ;
  wire \PCI-PAR/PER_4845 ;
  wire \PCI-PAR/P0I ;
  wire \PCI-PAR/X0I ;
  wire \PCI-PAR/X1I ;
  wire \PCI-PAR/P1I ;
  wire \PCI-PAR/X2I ;
  wire \PCI-PAR/X3I ;
  wire \PCI-PAR/P2I ;
  wire \PCI-PAR/X4I ;
  wire \PCI-PAR/X5I ;
  wire \PCI-PAR/P3I ;
  wire \PCI-PAR/X6I ;
  wire \PCI-PAR/X7I ;
  wire \PCI-PAR/$3I3033/$1N2216 ;
  wire \PCI-PAR/$3I3034/$1N2216 ;
  wire \PCI-PAR/$4I3135/$1N2216 ;
  wire \PCI-PAR/$4I3136/$1N2216 ;
  wire \PCI-PAR/$7I2990/$1N2216 ;
  wire \PCI-PAR/$7I2997/$1N2216 ;
  wire \$3I3124/$1N2216 ;
  wire \$3I3125/$1N2216 ;
  wire \$3I3126/$1N2216 ;
  wire \$3I3127/$1N2216 ;
  wire \$3I3128/$1N2216 ;
  wire \$3I3355/$1N2216 ;
  wire \$3I3356/$1N2216 ;
  wire \$3I3357/$1N2216 ;
  wire \$3I3358/$1N2216 ;
  wire \$3I3359/$1N2216 ;
  wire \BAR0/CSRENNL ;
  wire \BAR0/ENABLENL ;
  wire \BAR0/NL_CE ;
  wire \BAR0/$2N3280 ;
  wire \BAR0/$2N3273 ;
  wire \BAR0/NS_NL_MEM ;
  wire \BAR0/NS_HITNL ;
  wire \BAR0/UNALIGN ;
  wire \BAR0/$1N3458 ;
  wire \BAR0/CSREN64 ;
  wire \BAR0/ENABLE32 ;
  wire \BAR0/CSREN32 ;
  wire \BAR0/MATCH ;
  wire \BAR0/$1N3366 ;
  wire \BAR0/$1N3368 ;
  wire \BAR0/$1N3380 ;
  wire \BAR0/$1N3369 ;
  wire \BAR0/BR-31-24/$1N3111 ;
  wire \BAR0/BR-31-24/$1N3099 ;
  wire \BAR0/BR-31-24/$1N3110 ;
  wire \BAR0/BR-31-24/IN1 ;
  wire \BAR0/BR-31-24/IN3 ;
  wire \BAR0/BR-31-24/RAWQ3 ;
  wire \BAR0/BR-31-24/RAWQ2 ;
  wire \BAR0/BR-31-24/RAWQ1 ;
  wire \BAR0/BR-31-24/RAWQ0 ;
  wire \BAR0/BR-31-24/IN2 ;
  wire \BAR0/BR-31-24/EQ32_5482 ;
  wire \BAR0/BR-31-24/EQ3 ;
  wire \BAR0/BR-31-24/EQ2 ;
  wire \BAR0/BR-31-24/EQ10_5479 ;
  wire \BAR0/BR-31-24/EQ1 ;
  wire \BAR0/BR-31-24/EQ0 ;
  wire \BAR0/BR-31-24/IN0 ;
  wire \BAR0/BR-31-24/$1N2992 ;
  wire \BAR0/BR-31-24/$1N2911 ;
  wire \BAR0/BR-31-24/$1N2993 ;
  wire \BAR0/BR-31-24/EQ76_5472 ;
  wire \BAR0/BR-31-24/EQ4 ;
  wire \BAR0/BR-31-24/EQ6 ;
  wire \BAR0/BR-31-24/EQ54_5469 ;
  wire \BAR0/BR-31-24/IN4 ;
  wire \BAR0/BR-31-24/RAWQ7 ;
  wire \BAR0/BR-31-24/RAWQ4 ;
  wire \BAR0/BR-31-24/RAWQ5 ;
  wire \BAR0/BR-31-24/IN6 ;
  wire \BAR0/BR-31-24/RAWQ6 ;
  wire \BAR0/BR-31-24/EQ7 ;
  wire \BAR0/BR-31-24/IN7 ;
  wire \BAR0/BR-31-24/EQ5 ;
  wire \BAR0/BR-31-24/IN5 ;
  wire \BAR0/BR-31-24/$1N2910 ;
  wire \BAR0/BR-31-24/$1I2909/$1N2216 ;
  wire \BAR0/BR-31-24/$1I2990/$1N2216 ;
  wire \BAR0/BR-31-24/$1I3091/$1N2216 ;
  wire \BAR0/BR-31-24/$1I3096/$1N2216 ;
  wire \BAR0/BR-23-16/$1N3111 ;
  wire \BAR0/BR-23-16/$1N3099 ;
  wire \BAR0/BR-23-16/$1N3110 ;
  wire \BAR0/BR-23-16/IN1 ;
  wire \BAR0/BR-23-16/IN3 ;
  wire \BAR0/BR-23-16/RAWQ3 ;
  wire \BAR0/BR-23-16/RAWQ2 ;
  wire \BAR0/BR-23-16/RAWQ1 ;
  wire \BAR0/BR-23-16/RAWQ0 ;
  wire \BAR0/BR-23-16/IN2 ;
  wire \BAR0/BR-23-16/EQ32_5554 ;
  wire \BAR0/BR-23-16/EQ3 ;
  wire \BAR0/BR-23-16/EQ2 ;
  wire \BAR0/BR-23-16/EQ10_5551 ;
  wire \BAR0/BR-23-16/EQ1 ;
  wire \BAR0/BR-23-16/EQ0 ;
  wire \BAR0/BR-23-16/IN0 ;
  wire \BAR0/BR-23-16/$1N2992 ;
  wire \BAR0/BR-23-16/$1N2911 ;
  wire \BAR0/BR-23-16/$1N2993 ;
  wire \BAR0/BR-23-16/EQ76_5544 ;
  wire \BAR0/BR-23-16/EQ4 ;
  wire \BAR0/BR-23-16/EQ6 ;
  wire \BAR0/BR-23-16/EQ54_5541 ;
  wire \BAR0/BR-23-16/IN4 ;
  wire \BAR0/BR-23-16/RAWQ7 ;
  wire \BAR0/BR-23-16/RAWQ4 ;
  wire \BAR0/BR-23-16/RAWQ5 ;
  wire \BAR0/BR-23-16/IN6 ;
  wire \BAR0/BR-23-16/RAWQ6 ;
  wire \BAR0/BR-23-16/EQ7 ;
  wire \BAR0/BR-23-16/IN7 ;
  wire \BAR0/BR-23-16/EQ5 ;
  wire \BAR0/BR-23-16/IN5 ;
  wire \BAR0/BR-23-16/$1N2910 ;
  wire \BAR0/BR-23-16/$1I2909/$1N2216 ;
  wire \BAR0/BR-23-16/$1I2990/$1N2216 ;
  wire \BAR0/BR-23-16/$1I3091/$1N2216 ;
  wire \BAR0/BR-23-16/$1I3096/$1N2216 ;
  wire \BAR0/BR-15-8/$1N3111 ;
  wire \BAR0/BR-15-8/$1N3099 ;
  wire \BAR0/BR-15-8/$1N3110 ;
  wire \BAR0/BR-15-8/IN1 ;
  wire \BAR0/BR-15-8/IN3 ;
  wire \BAR0/BR-15-8/RAWQ3 ;
  wire \BAR0/BR-15-8/RAWQ2 ;
  wire \BAR0/BR-15-8/RAWQ1 ;
  wire \BAR0/BR-15-8/RAWQ0 ;
  wire \BAR0/BR-15-8/IN2 ;
  wire \BAR0/BR-15-8/EQ32_5626 ;
  wire \BAR0/BR-15-8/EQ3 ;
  wire \BAR0/BR-15-8/EQ2 ;
  wire \BAR0/BR-15-8/EQ10_5623 ;
  wire \BAR0/BR-15-8/EQ1 ;
  wire \BAR0/BR-15-8/EQ0 ;
  wire \BAR0/BR-15-8/IN0 ;
  wire \BAR0/BR-15-8/$1N2992 ;
  wire \BAR0/BR-15-8/$1N2911 ;
  wire \BAR0/BR-15-8/$1N2993 ;
  wire \BAR0/BR-15-8/EQ76_5616 ;
  wire \BAR0/BR-15-8/EQ4 ;
  wire \BAR0/BR-15-8/EQ6 ;
  wire \BAR0/BR-15-8/EQ54_5613 ;
  wire \BAR0/BR-15-8/IN4 ;
  wire \BAR0/BR-15-8/RAWQ7 ;
  wire \BAR0/BR-15-8/RAWQ4 ;
  wire \BAR0/BR-15-8/RAWQ5 ;
  wire \BAR0/BR-15-8/IN6 ;
  wire \BAR0/BR-15-8/RAWQ6 ;
  wire \BAR0/BR-15-8/EQ7 ;
  wire \BAR0/BR-15-8/IN7 ;
  wire \BAR0/BR-15-8/EQ5 ;
  wire \BAR0/BR-15-8/IN5 ;
  wire \BAR0/BR-15-8/$1N2910 ;
  wire \BAR0/BR-15-8/$1I2909/$1N2216 ;
  wire \BAR0/BR-15-8/$1I2990/$1N2216 ;
  wire \BAR0/BR-15-8/$1I3091/$1N2216 ;
  wire \BAR0/BR-15-8/$1I3096/$1N2216 ;
  wire \BAR0/BR-CMD/EX_N ;
  wire \BAR0/BR-CMD/MEM_5666 ;
  wire \BAR0/BR-CMD/$1N195 ;
  wire \BAR0/BR-CMD/$1N201 ;
  wire \BAR0/BR-CMD/IO_5663 ;
  wire \BAR0/BR-CMD/SEL ;
  wire \BAR0/BR-CMD/$1N144 ;
  wire \BAR0/BR-CMD/$1I143/$1N2216 ;
  wire \BAR0/BR-CMD/$1I223/M0 ;
  wire \BAR0/BR-CMD/$1I223/M1 ;
  wire \BAR0/BR-7-4/$1N2701 ;
  wire \BAR0/BR-7-4/$1N2706 ;
  wire \BAR0/BR-7-4/$1N2697 ;
  wire \BAR0/BR-7-4/EQ54_5702 ;
  wire \BAR0/BR-7-4/EQ76_5701 ;
  wire \BAR0/BR-7-4/EQ7 ;
  wire \BAR0/BR-7-4/IN7 ;
  wire \BAR0/BR-7-4/EQ6 ;
  wire \BAR0/BR-7-4/IN6 ;
  wire \BAR0/BR-7-4/EQ5 ;
  wire \BAR0/BR-7-4/IN5 ;
  wire \BAR0/BR-7-4/EQ4 ;
  wire \BAR0/BR-7-4/IN4 ;
  wire \BAR0/BR-7-4/RAWQ7 ;
  wire \BAR0/BR-7-4/RAWQ6 ;
  wire \BAR0/BR-7-4/RAWQ5 ;
  wire \BAR0/BR-7-4/RAWQ4 ;
  wire \BAR0/BR-7-4/$1I2700/$1N2216 ;
  wire \BAR0/BR-7-4/$1I2705/$1N2216 ;
  wire \BAR0/$1I3440/M0 ;
  wire \BAR0/$1I3440/M1 ;
  wire \BAR0/$1I3453/M0 ;
  wire \BAR0/$1I3453/M1 ;
  wire \BAR0/$1I3468/$1N2216 ;
  wire \BAR0/$1I3469/$1N2216 ;
  wire \BAR0/$2I3304/$1N2216 ;
  wire \BAR0/$2I3321/M0 ;
  wire \BAR0/$2I3321/M1 ;
  wire \BAR1/CSRENNL ;
  wire \BAR1/ENABLENL ;
  wire \BAR1/NL_CE ;
  wire \BAR1/$2N3280 ;
  wire \BAR1/$2N3273 ;
  wire \BAR1/NS_NL_MEM ;
  wire \BAR1/NS_HITNL ;
  wire \BAR1/UNALIGN ;
  wire \BAR1/$1N3458 ;
  wire \BAR1/CSREN64 ;
  wire \BAR1/ENABLE32 ;
  wire \BAR1/CSREN32 ;
  wire \BAR1/MATCH ;
  wire \BAR1/$1N3366 ;
  wire \BAR1/$1N3368 ;
  wire \BAR1/$1N3380 ;
  wire \BAR1/$1N3369 ;
  wire \BAR1/BR-31-24/$1N3111 ;
  wire \BAR1/BR-31-24/$1N3099 ;
  wire \BAR1/BR-31-24/$1N3110 ;
  wire \BAR1/BR-31-24/IN1 ;
  wire \BAR1/BR-31-24/IN3 ;
  wire \BAR1/BR-31-24/RAWQ3 ;
  wire \BAR1/BR-31-24/RAWQ2 ;
  wire \BAR1/BR-31-24/RAWQ1 ;
  wire \BAR1/BR-31-24/RAWQ0 ;
  wire \BAR1/BR-31-24/IN2 ;
  wire \BAR1/BR-31-24/EQ32_5941 ;
  wire \BAR1/BR-31-24/EQ3 ;
  wire \BAR1/BR-31-24/EQ2 ;
  wire \BAR1/BR-31-24/EQ10_5938 ;
  wire \BAR1/BR-31-24/EQ1 ;
  wire \BAR1/BR-31-24/EQ0 ;
  wire \BAR1/BR-31-24/IN0 ;
  wire \BAR1/BR-31-24/$1N2992 ;
  wire \BAR1/BR-31-24/$1N2911 ;
  wire \BAR1/BR-31-24/$1N2993 ;
  wire \BAR1/BR-31-24/EQ76_5931 ;
  wire \BAR1/BR-31-24/EQ4 ;
  wire \BAR1/BR-31-24/EQ6 ;
  wire \BAR1/BR-31-24/EQ54_5928 ;
  wire \BAR1/BR-31-24/IN4 ;
  wire \BAR1/BR-31-24/RAWQ7 ;
  wire \BAR1/BR-31-24/RAWQ4 ;
  wire \BAR1/BR-31-24/RAWQ5 ;
  wire \BAR1/BR-31-24/IN6 ;
  wire \BAR1/BR-31-24/RAWQ6 ;
  wire \BAR1/BR-31-24/EQ7 ;
  wire \BAR1/BR-31-24/IN7 ;
  wire \BAR1/BR-31-24/EQ5 ;
  wire \BAR1/BR-31-24/IN5 ;
  wire \BAR1/BR-31-24/$1N2910 ;
  wire \BAR1/BR-31-24/$1I2909/$1N2216 ;
  wire \BAR1/BR-31-24/$1I2990/$1N2216 ;
  wire \BAR1/BR-31-24/$1I3091/$1N2216 ;
  wire \BAR1/BR-31-24/$1I3096/$1N2216 ;
  wire \BAR1/BR-23-16/$1N3111 ;
  wire \BAR1/BR-23-16/$1N3099 ;
  wire \BAR1/BR-23-16/$1N3110 ;
  wire \BAR1/BR-23-16/IN1 ;
  wire \BAR1/BR-23-16/IN3 ;
  wire \BAR1/BR-23-16/RAWQ3 ;
  wire \BAR1/BR-23-16/RAWQ2 ;
  wire \BAR1/BR-23-16/RAWQ1 ;
  wire \BAR1/BR-23-16/RAWQ0 ;
  wire \BAR1/BR-23-16/IN2 ;
  wire \BAR1/BR-23-16/EQ32_6013 ;
  wire \BAR1/BR-23-16/EQ3 ;
  wire \BAR1/BR-23-16/EQ2 ;
  wire \BAR1/BR-23-16/EQ10_6010 ;
  wire \BAR1/BR-23-16/EQ1 ;
  wire \BAR1/BR-23-16/EQ0 ;
  wire \BAR1/BR-23-16/IN0 ;
  wire \BAR1/BR-23-16/$1N2992 ;
  wire \BAR1/BR-23-16/$1N2911 ;
  wire \BAR1/BR-23-16/$1N2993 ;
  wire \BAR1/BR-23-16/EQ76_6003 ;
  wire \BAR1/BR-23-16/EQ4 ;
  wire \BAR1/BR-23-16/EQ6 ;
  wire \BAR1/BR-23-16/EQ54_6000 ;
  wire \BAR1/BR-23-16/IN4 ;
  wire \BAR1/BR-23-16/RAWQ7 ;
  wire \BAR1/BR-23-16/RAWQ4 ;
  wire \BAR1/BR-23-16/RAWQ5 ;
  wire \BAR1/BR-23-16/IN6 ;
  wire \BAR1/BR-23-16/RAWQ6 ;
  wire \BAR1/BR-23-16/EQ7 ;
  wire \BAR1/BR-23-16/IN7 ;
  wire \BAR1/BR-23-16/EQ5 ;
  wire \BAR1/BR-23-16/IN5 ;
  wire \BAR1/BR-23-16/$1N2910 ;
  wire \BAR1/BR-23-16/$1I2909/$1N2216 ;
  wire \BAR1/BR-23-16/$1I2990/$1N2216 ;
  wire \BAR1/BR-23-16/$1I3091/$1N2216 ;
  wire \BAR1/BR-23-16/$1I3096/$1N2216 ;
  wire \BAR1/BR-15-8/$1N3111 ;
  wire \BAR1/BR-15-8/$1N3099 ;
  wire \BAR1/BR-15-8/$1N3110 ;
  wire \BAR1/BR-15-8/IN1 ;
  wire \BAR1/BR-15-8/IN3 ;
  wire \BAR1/BR-15-8/RAWQ3 ;
  wire \BAR1/BR-15-8/RAWQ2 ;
  wire \BAR1/BR-15-8/RAWQ1 ;
  wire \BAR1/BR-15-8/RAWQ0 ;
  wire \BAR1/BR-15-8/IN2 ;
  wire \BAR1/BR-15-8/EQ32_6085 ;
  wire \BAR1/BR-15-8/EQ3 ;
  wire \BAR1/BR-15-8/EQ2 ;
  wire \BAR1/BR-15-8/EQ10_6082 ;
  wire \BAR1/BR-15-8/EQ1 ;
  wire \BAR1/BR-15-8/EQ0 ;
  wire \BAR1/BR-15-8/IN0 ;
  wire \BAR1/BR-15-8/$1N2992 ;
  wire \BAR1/BR-15-8/$1N2911 ;
  wire \BAR1/BR-15-8/$1N2993 ;
  wire \BAR1/BR-15-8/EQ76_6075 ;
  wire \BAR1/BR-15-8/EQ4 ;
  wire \BAR1/BR-15-8/EQ6 ;
  wire \BAR1/BR-15-8/EQ54_6072 ;
  wire \BAR1/BR-15-8/IN4 ;
  wire \BAR1/BR-15-8/RAWQ7 ;
  wire \BAR1/BR-15-8/RAWQ4 ;
  wire \BAR1/BR-15-8/RAWQ5 ;
  wire \BAR1/BR-15-8/IN6 ;
  wire \BAR1/BR-15-8/RAWQ6 ;
  wire \BAR1/BR-15-8/EQ7 ;
  wire \BAR1/BR-15-8/IN7 ;
  wire \BAR1/BR-15-8/EQ5 ;
  wire \BAR1/BR-15-8/IN5 ;
  wire \BAR1/BR-15-8/$1N2910 ;
  wire \BAR1/BR-15-8/$1I2909/$1N2216 ;
  wire \BAR1/BR-15-8/$1I2990/$1N2216 ;
  wire \BAR1/BR-15-8/$1I3091/$1N2216 ;
  wire \BAR1/BR-15-8/$1I3096/$1N2216 ;
  wire \BAR1/BR-CMD/EX_N ;
  wire \BAR1/BR-CMD/MEM_6125 ;
  wire \BAR1/BR-CMD/$1N195 ;
  wire \BAR1/BR-CMD/$1N201 ;
  wire \BAR1/BR-CMD/IO_6122 ;
  wire \BAR1/BR-CMD/SEL ;
  wire \BAR1/BR-CMD/$1N144 ;
  wire \BAR1/BR-CMD/$1I143/$1N2216 ;
  wire \BAR1/BR-CMD/$1I223/M0 ;
  wire \BAR1/BR-CMD/$1I223/M1 ;
  wire \BAR1/BR-7-4/$1N2701 ;
  wire \BAR1/BR-7-4/$1N2706 ;
  wire \BAR1/BR-7-4/$1N2697 ;
  wire \BAR1/BR-7-4/EQ54_6161 ;
  wire \BAR1/BR-7-4/EQ76_6160 ;
  wire \BAR1/BR-7-4/EQ7 ;
  wire \BAR1/BR-7-4/IN7 ;
  wire \BAR1/BR-7-4/EQ6 ;
  wire \BAR1/BR-7-4/IN6 ;
  wire \BAR1/BR-7-4/EQ5 ;
  wire \BAR1/BR-7-4/IN5 ;
  wire \BAR1/BR-7-4/EQ4 ;
  wire \BAR1/BR-7-4/IN4 ;
  wire \BAR1/BR-7-4/RAWQ7 ;
  wire \BAR1/BR-7-4/RAWQ6 ;
  wire \BAR1/BR-7-4/RAWQ5 ;
  wire \BAR1/BR-7-4/RAWQ4 ;
  wire \BAR1/BR-7-4/$1I2700/$1N2216 ;
  wire \BAR1/BR-7-4/$1I2705/$1N2216 ;
  wire \BAR1/$1I3440/M0 ;
  wire \BAR1/$1I3440/M1 ;
  wire \BAR1/$1I3453/M0 ;
  wire \BAR1/$1I3453/M1 ;
  wire \BAR1/$1I3468/$1N2216 ;
  wire \BAR1/$1I3469/$1N2216 ;
  wire \BAR1/$2I3304/$1N2216 ;
  wire \BAR1/$2I3321/M0 ;
  wire \BAR1/$2I3321/M1 ;
  wire \BAR2/CSRENNL ;
  wire \BAR2/ENABLENL ;
  wire \BAR2/NL_CE ;
  wire \BAR2/$2N3280 ;
  wire \BAR2/$2N3273 ;
  wire \BAR2/NS_NL_MEM ;
  wire \BAR2/NS_HITNL ;
  wire \BAR2/UNALIGN ;
  wire \BAR2/$1N3458 ;
  wire \BAR2/CSREN64 ;
  wire \BAR2/ENABLE32 ;
  wire \BAR2/CSREN32 ;
  wire \BAR2/MATCH ;
  wire \BAR2/$1N3366 ;
  wire \BAR2/$1N3368 ;
  wire \BAR2/$1N3380 ;
  wire \BAR2/$1N3369 ;
  wire \BAR2/BR-31-24/$1N3111 ;
  wire \BAR2/BR-31-24/$1N3099 ;
  wire \BAR2/BR-31-24/$1N3110 ;
  wire \BAR2/BR-31-24/IN1 ;
  wire \BAR2/BR-31-24/IN3 ;
  wire \BAR2/BR-31-24/RAWQ3 ;
  wire \BAR2/BR-31-24/RAWQ2 ;
  wire \BAR2/BR-31-24/RAWQ1 ;
  wire \BAR2/BR-31-24/RAWQ0 ;
  wire \BAR2/BR-31-24/IN2 ;
  wire \BAR2/BR-31-24/EQ32_6400 ;
  wire \BAR2/BR-31-24/EQ3 ;
  wire \BAR2/BR-31-24/EQ2 ;
  wire \BAR2/BR-31-24/EQ10_6397 ;
  wire \BAR2/BR-31-24/EQ1 ;
  wire \BAR2/BR-31-24/EQ0 ;
  wire \BAR2/BR-31-24/IN0 ;
  wire \BAR2/BR-31-24/$1N2992 ;
  wire \BAR2/BR-31-24/$1N2911 ;
  wire \BAR2/BR-31-24/$1N2993 ;
  wire \BAR2/BR-31-24/EQ76_6390 ;
  wire \BAR2/BR-31-24/EQ4 ;
  wire \BAR2/BR-31-24/EQ6 ;
  wire \BAR2/BR-31-24/EQ54_6387 ;
  wire \BAR2/BR-31-24/IN4 ;
  wire \BAR2/BR-31-24/RAWQ7 ;
  wire \BAR2/BR-31-24/RAWQ4 ;
  wire \BAR2/BR-31-24/RAWQ5 ;
  wire \BAR2/BR-31-24/IN6 ;
  wire \BAR2/BR-31-24/RAWQ6 ;
  wire \BAR2/BR-31-24/EQ7 ;
  wire \BAR2/BR-31-24/IN7 ;
  wire \BAR2/BR-31-24/EQ5 ;
  wire \BAR2/BR-31-24/IN5 ;
  wire \BAR2/BR-31-24/$1N2910 ;
  wire \BAR2/BR-31-24/$1I2909/$1N2216 ;
  wire \BAR2/BR-31-24/$1I2990/$1N2216 ;
  wire \BAR2/BR-31-24/$1I3091/$1N2216 ;
  wire \BAR2/BR-31-24/$1I3096/$1N2216 ;
  wire \BAR2/BR-23-16/$1N3111 ;
  wire \BAR2/BR-23-16/$1N3099 ;
  wire \BAR2/BR-23-16/$1N3110 ;
  wire \BAR2/BR-23-16/IN1 ;
  wire \BAR2/BR-23-16/IN3 ;
  wire \BAR2/BR-23-16/RAWQ3 ;
  wire \BAR2/BR-23-16/RAWQ2 ;
  wire \BAR2/BR-23-16/RAWQ1 ;
  wire \BAR2/BR-23-16/RAWQ0 ;
  wire \BAR2/BR-23-16/IN2 ;
  wire \BAR2/BR-23-16/EQ32_6472 ;
  wire \BAR2/BR-23-16/EQ3 ;
  wire \BAR2/BR-23-16/EQ2 ;
  wire \BAR2/BR-23-16/EQ10_6469 ;
  wire \BAR2/BR-23-16/EQ1 ;
  wire \BAR2/BR-23-16/EQ0 ;
  wire \BAR2/BR-23-16/IN0 ;
  wire \BAR2/BR-23-16/$1N2992 ;
  wire \BAR2/BR-23-16/$1N2911 ;
  wire \BAR2/BR-23-16/$1N2993 ;
  wire \BAR2/BR-23-16/EQ76_6462 ;
  wire \BAR2/BR-23-16/EQ4 ;
  wire \BAR2/BR-23-16/EQ6 ;
  wire \BAR2/BR-23-16/EQ54_6459 ;
  wire \BAR2/BR-23-16/IN4 ;
  wire \BAR2/BR-23-16/RAWQ7 ;
  wire \BAR2/BR-23-16/RAWQ4 ;
  wire \BAR2/BR-23-16/RAWQ5 ;
  wire \BAR2/BR-23-16/IN6 ;
  wire \BAR2/BR-23-16/RAWQ6 ;
  wire \BAR2/BR-23-16/EQ7 ;
  wire \BAR2/BR-23-16/IN7 ;
  wire \BAR2/BR-23-16/EQ5 ;
  wire \BAR2/BR-23-16/IN5 ;
  wire \BAR2/BR-23-16/$1N2910 ;
  wire \BAR2/BR-23-16/$1I2909/$1N2216 ;
  wire \BAR2/BR-23-16/$1I2990/$1N2216 ;
  wire \BAR2/BR-23-16/$1I3091/$1N2216 ;
  wire \BAR2/BR-23-16/$1I3096/$1N2216 ;
  wire \BAR2/BR-15-8/$1N3111 ;
  wire \BAR2/BR-15-8/$1N3099 ;
  wire \BAR2/BR-15-8/$1N3110 ;
  wire \BAR2/BR-15-8/IN1 ;
  wire \BAR2/BR-15-8/IN3 ;
  wire \BAR2/BR-15-8/RAWQ3 ;
  wire \BAR2/BR-15-8/RAWQ2 ;
  wire \BAR2/BR-15-8/RAWQ1 ;
  wire \BAR2/BR-15-8/RAWQ0 ;
  wire \BAR2/BR-15-8/IN2 ;
  wire \BAR2/BR-15-8/EQ32_6544 ;
  wire \BAR2/BR-15-8/EQ3 ;
  wire \BAR2/BR-15-8/EQ2 ;
  wire \BAR2/BR-15-8/EQ10_6541 ;
  wire \BAR2/BR-15-8/EQ1 ;
  wire \BAR2/BR-15-8/EQ0 ;
  wire \BAR2/BR-15-8/IN0 ;
  wire \BAR2/BR-15-8/$1N2992 ;
  wire \BAR2/BR-15-8/$1N2911 ;
  wire \BAR2/BR-15-8/$1N2993 ;
  wire \BAR2/BR-15-8/EQ76_6534 ;
  wire \BAR2/BR-15-8/EQ4 ;
  wire \BAR2/BR-15-8/EQ6 ;
  wire \BAR2/BR-15-8/EQ54_6531 ;
  wire \BAR2/BR-15-8/IN4 ;
  wire \BAR2/BR-15-8/RAWQ7 ;
  wire \BAR2/BR-15-8/RAWQ4 ;
  wire \BAR2/BR-15-8/RAWQ5 ;
  wire \BAR2/BR-15-8/IN6 ;
  wire \BAR2/BR-15-8/RAWQ6 ;
  wire \BAR2/BR-15-8/EQ7 ;
  wire \BAR2/BR-15-8/IN7 ;
  wire \BAR2/BR-15-8/EQ5 ;
  wire \BAR2/BR-15-8/IN5 ;
  wire \BAR2/BR-15-8/$1N2910 ;
  wire \BAR2/BR-15-8/$1I2909/$1N2216 ;
  wire \BAR2/BR-15-8/$1I2990/$1N2216 ;
  wire \BAR2/BR-15-8/$1I3091/$1N2216 ;
  wire \BAR2/BR-15-8/$1I3096/$1N2216 ;
  wire \BAR2/BR-CMD/EX_N ;
  wire \BAR2/BR-CMD/MEM_6584 ;
  wire \BAR2/BR-CMD/$1N195 ;
  wire \BAR2/BR-CMD/$1N201 ;
  wire \BAR2/BR-CMD/IO_6581 ;
  wire \BAR2/BR-CMD/SEL ;
  wire \BAR2/BR-CMD/$1N144 ;
  wire \BAR2/BR-CMD/$1I143/$1N2216 ;
  wire \BAR2/BR-CMD/$1I223/M0 ;
  wire \BAR2/BR-CMD/$1I223/M1 ;
  wire \BAR2/BR-7-4/$1N2701 ;
  wire \BAR2/BR-7-4/$1N2706 ;
  wire \BAR2/BR-7-4/$1N2697 ;
  wire \BAR2/BR-7-4/EQ54_6620 ;
  wire \BAR2/BR-7-4/EQ76_6619 ;
  wire \BAR2/BR-7-4/EQ7 ;
  wire \BAR2/BR-7-4/IN7 ;
  wire \BAR2/BR-7-4/EQ6 ;
  wire \BAR2/BR-7-4/IN6 ;
  wire \BAR2/BR-7-4/EQ5 ;
  wire \BAR2/BR-7-4/IN5 ;
  wire \BAR2/BR-7-4/EQ4 ;
  wire \BAR2/BR-7-4/IN4 ;
  wire \BAR2/BR-7-4/RAWQ7 ;
  wire \BAR2/BR-7-4/RAWQ6 ;
  wire \BAR2/BR-7-4/RAWQ5 ;
  wire \BAR2/BR-7-4/RAWQ4 ;
  wire \BAR2/BR-7-4/$1I2700/$1N2216 ;
  wire \BAR2/BR-7-4/$1I2705/$1N2216 ;
  wire \BAR2/$1I3440/M0 ;
  wire \BAR2/$1I3440/M1 ;
  wire \BAR2/$1I3453/M0 ;
  wire \BAR2/$1I3453/M1 ;
  wire \BAR2/$1I3468/$1N2216 ;
  wire \BAR2/$1I3469/$1N2216 ;
  wire \BAR2/$2I3304/$1N2216 ;
  wire \BAR2/$2I3321/M0 ;
  wire \BAR2/$2I3321/M1 ;
  wire \PCI-IREG/INT-PINX/$1I2486/$1N2216 ;
  wire \PCI-IREG/INT-PINX/$1I2488/$1N2216 ;
  wire \PCI-IREG/INT-PINX/$1I2490/$1N2216 ;
  wire \PCI-IREG/INT-PINX/$1I2492/$1N2216 ;
  wire \PCI-IREG/INT-PINX/$1I2494/$1N2216 ;
  wire \PCI-IREG/INT-PINX/$1I2496/$1N2216 ;
  wire \PCI-IREG/INT-PINX/$1I2498/$1N2216 ;
  wire \PCI-CSR/CMDREG/$1N2560 ;
  wire \PCI-CSR/CMDREG/$1N2556 ;
  wire \PCI-CSR/CMDREG/$1N2562 ;
  wire \PCI-CSR/CMDREG/$1N2559 ;
  wire \PCI-CSR/CMDREG/$1N2514 ;
  wire \PCI-CSR/CMDREG/$1N2527 ;
  wire \PCI-CSR/CMDREG/$1N2524 ;
  wire \PCI-CSR/CMDREG/$1N2525 ;
  wire \PCI-CSR/CMDREG/$1N2523 ;
  wire \PCI-CSR/CMDREG/$1N2522 ;
  wire \PCI-CSR/CMDREG/$1N2446 ;
  wire \PCI-CSR/CMDREG/$1N2346 ;
  wire \PCI-CSR/CMDREG/$1I2520/$1N2216 ;
  wire \PCI-CSR/CMDREG/$1I2521/$1N2216 ;
  wire \PCI-CSR/CMDREG/$1I2528/$1N2216 ;
  wire \PCI-CSR/CMDREG/$1I2529/$1N2216 ;
  wire \PCI-CSR/CMDREG/$1I2530/$1N2216 ;
  wire \PCI-CSR/CMDREG/$1I2532/$1N2216 ;
  wire \PCI-CSR/CMDREG/$1I2557/$1N2216 ;
  wire \PCI-CSR/CMDREG/$1I2558/$1N2216 ;
  wire \PCI-CSR/CMDREG/$1I2561/$1N2216 ;
  wire \PCI-CSR/CMDREG/$1I2583/$1N2216 ;
  wire \PCI-CSR/STATREG/$1N2634 ;
  wire \PCI-CSR/STATREG/$1N2630 ;
  wire \PCI-CSR/STATREG/$1N2595 ;
  wire \PCI-CSR/STATREG/$1N2588 ;
  wire \PCI-CSR/STATREG/$1N2585 ;
  wire \PCI-CSR/STATREG/$1N2474 ;
  wire \PCI-CSR/STATREG/$1N2605 ;
  wire \PCI-CSR/STATREG/$1N2606 ;
  wire \PCI-CSR/STATREG/$1N2609 ;
  wire \PCI-CSR/STATREG/Q14/$1N2238 ;
  wire \PCI-CSR/STATREG/Q14/$1N2240 ;
  wire \PCI-CSR/STATREG/Q14/D ;
  wire \PCI-CSR/STATREG/Q14/$1I2233/M1 ;
  wire \PCI-CSR/STATREG/Q14/$1I2233/M0 ;
  wire \PCI-CSR/STATREG/Q12/$1N2238 ;
  wire \PCI-CSR/STATREG/Q12/$1N2240 ;
  wire \PCI-CSR/STATREG/Q12/D ;
  wire \PCI-CSR/STATREG/Q12/$1I2233/M1 ;
  wire \PCI-CSR/STATREG/Q12/$1I2233/M0 ;
  wire \PCI-CSR/STATREG/Q8/$1N2238 ;
  wire \PCI-CSR/STATREG/Q8/$1N2240 ;
  wire \PCI-CSR/STATREG/Q8/D ;
  wire \PCI-CSR/STATREG/Q8/$1I2233/M1 ;
  wire \PCI-CSR/STATREG/Q8/$1I2233/M0 ;
  wire \PCI-CSR/STATREG/Q11/$1N2238 ;
  wire \PCI-CSR/STATREG/Q11/$1N2240 ;
  wire \PCI-CSR/STATREG/Q11/D ;
  wire \PCI-CSR/STATREG/Q11/$1I2233/M1 ;
  wire \PCI-CSR/STATREG/Q11/$1I2233/M0 ;
  wire \PCI-CSR/STATREG/Q13/$1N2238 ;
  wire \PCI-CSR/STATREG/Q13/$1N2240 ;
  wire \PCI-CSR/STATREG/Q13/D ;
  wire \PCI-CSR/STATREG/Q13/$1I2233/M1 ;
  wire \PCI-CSR/STATREG/Q13/$1I2233/M0 ;
  wire \PCI-CSR/STATREG/Q15/$1N2238 ;
  wire \PCI-CSR/STATREG/Q15/$1N2240 ;
  wire \PCI-CSR/STATREG/Q15/D ;
  wire \PCI-CSR/STATREG/Q15/$1I2233/M1 ;
  wire \PCI-CSR/STATREG/Q15/$1I2233/M0 ;
  wire \PCI-CSR/STATREG/$1I2569/$1N2216 ;
  wire \PCI-CSR/STATREG/$1I2587/$1N2216 ;
  wire \PCI-CSR/STATREG/$1I2590/$1N2216 ;
  wire \PCI-CSR/STATREG/$1I2596/$1N2216 ;
  wire \PCI-CSR/STATREG/$1I2604/$1N2216 ;
  wire \PCI-CSR/STATREG/$1I2607/$1N2216 ;
  wire \PCI-CSR/STATREG/$1I2608/$1N2216 ;
  wire \PCI-CSR/STATREG/$1I2631/$1N2216 ;
  wire \PCI-ROM/ROM0 ;
  wire \PCI-ROM/ROM1 ;
  wire \PCI-ROM/ROM2 ;
  wire \PCI-ROM/ROM3 ;
  wire \PCI-ROM/ROM4 ;
  wire \PCI-ROM/ROM5 ;
  wire \PCI-ROM/ROM6 ;
  wire \PCI-ROM/ROM7 ;
  wire \PCI-ROM/ROM8 ;
  wire \PCI-ROM/ROM9 ;
  wire \PCI-ROM/ROM10 ;
  wire \PCI-ROM/ROM11 ;
  wire \PCI-ROM/ROM12 ;
  wire \PCI-ROM/ROM13 ;
  wire \PCI-ROM/ROM14 ;
  wire \PCI-ROM/ROM15 ;
  wire \PCI-ROM/ROM16 ;
  wire \PCI-ROM/ROM17 ;
  wire \PCI-ROM/ROM18 ;
  wire \PCI-ROM/ROM19 ;
  wire \PCI-ROM/ROM20 ;
  wire \PCI-ROM/ROM21 ;
  wire \PCI-ROM/ROM22 ;
  wire \PCI-ROM/ROM23 ;
  wire \PCI-ROM/ROM24 ;
  wire \PCI-ROM/ROM25 ;
  wire \PCI-ROM/ROM26 ;
  wire \PCI-ROM/ROM27 ;
  wire \PCI-ROM/ROM28 ;
  wire \PCI-ROM/ROM29 ;
  wire \PCI-ROM/ROM30 ;
  wire \PCI-ROM/ROM31 ;
  wire \PCI-ROM/$1N8453 ;
  wire \PCI-ROM/RF0 ;
  wire \PCI-ROM/CLR0 ;
  wire \PCI-ROM/RF1 ;
  wire \PCI-ROM/CLR1 ;
  wire \PCI-ROM/RF2 ;
  wire \PCI-ROM/CLR2 ;
  wire \PCI-ROM/RF3 ;
  wire \PCI-ROM/CLR3 ;
  wire \PCI-ROM/RF4 ;
  wire \PCI-ROM/CLR4 ;
  wire \PCI-ROM/RF5 ;
  wire \PCI-ROM/CLR5 ;
  wire \PCI-ROM/RF6 ;
  wire \PCI-ROM/CLR6 ;
  wire \PCI-ROM/RF7 ;
  wire \PCI-ROM/CLR7 ;
  wire \PCI-ROM/RF8 ;
  wire \PCI-ROM/CLR8 ;
  wire \PCI-ROM/RF9 ;
  wire \PCI-ROM/CLR9 ;
  wire \PCI-ROM/RF10 ;
  wire \PCI-ROM/CLR10 ;
  wire \PCI-ROM/RF11 ;
  wire \PCI-ROM/CLR11 ;
  wire \PCI-ROM/RF12 ;
  wire \PCI-ROM/CLR12 ;
  wire \PCI-ROM/RF13 ;
  wire \PCI-ROM/CLR13 ;
  wire \PCI-ROM/RF14 ;
  wire \PCI-ROM/CLR14 ;
  wire \PCI-ROM/RF15 ;
  wire \PCI-ROM/CLR15 ;
  wire \PCI-ROM/RF16 ;
  wire \PCI-ROM/CLR16 ;
  wire \PCI-ROM/RF17 ;
  wire \PCI-ROM/CLR17 ;
  wire \PCI-ROM/RF18 ;
  wire \PCI-ROM/CLR18 ;
  wire \PCI-ROM/RF19 ;
  wire \PCI-ROM/CLR19 ;
  wire \PCI-ROM/RF20 ;
  wire \PCI-ROM/CLR20 ;
  wire \PCI-ROM/RF21 ;
  wire \PCI-ROM/CLR21 ;
  wire \PCI-ROM/RF22 ;
  wire \PCI-ROM/CLR22 ;
  wire \PCI-ROM/RF23 ;
  wire \PCI-ROM/CLR23 ;
  wire \PCI-ROM/RF24 ;
  wire \PCI-ROM/CLR24 ;
  wire \PCI-ROM/RF25 ;
  wire \PCI-ROM/CLR25 ;
  wire \PCI-ROM/RF26 ;
  wire \PCI-ROM/CLR26 ;
  wire \PCI-ROM/RF27 ;
  wire \PCI-ROM/CLR27 ;
  wire \PCI-ROM/RF28 ;
  wire \PCI-ROM/CLR28 ;
  wire \PCI-ROM/RF29 ;
  wire \PCI-ROM/CLR29 ;
  wire \PCI-ROM/RF30 ;
  wire \PCI-ROM/CLR30 ;
  wire \PCI-ROM/RF31 ;
  wire \PCI-ROM/CLR31 ;
  wire \PCI-ROM/SELD ;
  wire \PCI-ROM/$1N8328 ;
  wire \PCI-ROM/RE0 ;
  wire \PCI-ROM/RE1 ;
  wire \PCI-ROM/RE2 ;
  wire \PCI-ROM/RE3 ;
  wire \PCI-ROM/RE4 ;
  wire \PCI-ROM/RE5 ;
  wire \PCI-ROM/RE6 ;
  wire \PCI-ROM/RE7 ;
  wire \PCI-ROM/RE8 ;
  wire \PCI-ROM/RE9 ;
  wire \PCI-ROM/RE10 ;
  wire \PCI-ROM/RE11 ;
  wire \PCI-ROM/RE12 ;
  wire \PCI-ROM/RE13 ;
  wire \PCI-ROM/RE14 ;
  wire \PCI-ROM/RE15 ;
  wire \PCI-ROM/RE16 ;
  wire \PCI-ROM/RE17 ;
  wire \PCI-ROM/RE18 ;
  wire \PCI-ROM/RE19 ;
  wire \PCI-ROM/RE20 ;
  wire \PCI-ROM/RE21 ;
  wire \PCI-ROM/RE22 ;
  wire \PCI-ROM/RE23 ;
  wire \PCI-ROM/RE24 ;
  wire \PCI-ROM/RE25 ;
  wire \PCI-ROM/RE26 ;
  wire \PCI-ROM/RE27 ;
  wire \PCI-ROM/RE28 ;
  wire \PCI-ROM/RE29 ;
  wire \PCI-ROM/RE30 ;
  wire \PCI-ROM/RE31 ;
  wire \PCI-ROM/SELBY ;
  wire \PCI-ROM/$1N8283 ;
  wire \PCI-ROM/RD0 ;
  wire \PCI-ROM/RD1 ;
  wire \PCI-ROM/RD2 ;
  wire \PCI-ROM/RD3 ;
  wire \PCI-ROM/RD4 ;
  wire \PCI-ROM/RD5 ;
  wire \PCI-ROM/RD6 ;
  wire \PCI-ROM/RD7 ;
  wire \PCI-ROM/RD8 ;
  wire \PCI-ROM/RD9 ;
  wire \PCI-ROM/RD10 ;
  wire \PCI-ROM/RD11 ;
  wire \PCI-ROM/RD12 ;
  wire \PCI-ROM/RD13 ;
  wire \PCI-ROM/RD14 ;
  wire \PCI-ROM/RD15 ;
  wire \PCI-ROM/RD16 ;
  wire \PCI-ROM/RD17 ;
  wire \PCI-ROM/RD18 ;
  wire \PCI-ROM/RD19 ;
  wire \PCI-ROM/RD20 ;
  wire \PCI-ROM/RD21 ;
  wire \PCI-ROM/RD22 ;
  wire \PCI-ROM/RD23 ;
  wire \PCI-ROM/RD24 ;
  wire \PCI-ROM/RD25 ;
  wire \PCI-ROM/RD26 ;
  wire \PCI-ROM/RD27 ;
  wire \PCI-ROM/RD28 ;
  wire \PCI-ROM/RD29 ;
  wire \PCI-ROM/RD30 ;
  wire \PCI-ROM/RD31 ;
  wire \PCI-ROM/SELBX ;
  wire \PCI-ROM/$1N8238 ;
  wire \PCI-ROM/$1N8188 ;
  wire \PCI-ROM/RC0 ;
  wire \PCI-ROM/RC1 ;
  wire \PCI-ROM/RC2 ;
  wire \PCI-ROM/RC3 ;
  wire \PCI-ROM/RC4 ;
  wire \PCI-ROM/RC5 ;
  wire \PCI-ROM/RC6 ;
  wire \PCI-ROM/RC7 ;
  wire \PCI-ROM/RC8 ;
  wire \PCI-ROM/RC9 ;
  wire \PCI-ROM/RC10 ;
  wire \PCI-ROM/RC11 ;
  wire \PCI-ROM/RC12 ;
  wire \PCI-ROM/RC13 ;
  wire \PCI-ROM/RC14 ;
  wire \PCI-ROM/RC15 ;
  wire \PCI-ROM/RC16 ;
  wire \PCI-ROM/RC17 ;
  wire \PCI-ROM/RC18 ;
  wire \PCI-ROM/RC19 ;
  wire \PCI-ROM/RC20 ;
  wire \PCI-ROM/RC21 ;
  wire \PCI-ROM/RC22 ;
  wire \PCI-ROM/RC23 ;
  wire \PCI-ROM/RC24 ;
  wire \PCI-ROM/RC25 ;
  wire \PCI-ROM/RC26 ;
  wire \PCI-ROM/RC27 ;
  wire \PCI-ROM/RC28 ;
  wire \PCI-ROM/RC29 ;
  wire \PCI-ROM/RC30 ;
  wire \PCI-ROM/RC31 ;
  wire \PCI-ROM/SELA ;
  wire \PCI-ROM/RA0 ;
  wire \PCI-ROM/RA1 ;
  wire \PCI-ROM/RA2 ;
  wire \PCI-ROM/RA3 ;
  wire \PCI-ROM/RA4 ;
  wire \PCI-ROM/RA5 ;
  wire \PCI-ROM/RA6 ;
  wire \PCI-ROM/RA7 ;
  wire \PCI-ROM/RA8 ;
  wire \PCI-ROM/RA9 ;
  wire \PCI-ROM/RA10 ;
  wire \PCI-ROM/RA11 ;
  wire \PCI-ROM/RA12 ;
  wire \PCI-ROM/RA13 ;
  wire \PCI-ROM/RA14 ;
  wire \PCI-ROM/RA15 ;
  wire \PCI-ROM/RA16 ;
  wire \PCI-ROM/RA17 ;
  wire \PCI-ROM/RA18 ;
  wire \PCI-ROM/RA19 ;
  wire \PCI-ROM/RA20 ;
  wire \PCI-ROM/RA21 ;
  wire \PCI-ROM/RA22 ;
  wire \PCI-ROM/RA23 ;
  wire \PCI-ROM/RA24 ;
  wire \PCI-ROM/RA25 ;
  wire \PCI-ROM/RA26 ;
  wire \PCI-ROM/RA27 ;
  wire \PCI-ROM/RA28 ;
  wire \PCI-ROM/RA29 ;
  wire \PCI-ROM/RA30 ;
  wire \PCI-ROM/RA31 ;
  wire \PCI-ROM/RB0 ;
  wire \PCI-ROM/RB1 ;
  wire \PCI-ROM/RB2 ;
  wire \PCI-ROM/RB3 ;
  wire \PCI-ROM/RB4 ;
  wire \PCI-ROM/RB5 ;
  wire \PCI-ROM/RB6 ;
  wire \PCI-ROM/RB7 ;
  wire \PCI-ROM/RB8 ;
  wire \PCI-ROM/RB9 ;
  wire \PCI-ROM/RB10 ;
  wire \PCI-ROM/RB11 ;
  wire \PCI-ROM/RB12 ;
  wire \PCI-ROM/RB13 ;
  wire \PCI-ROM/RB14 ;
  wire \PCI-ROM/RB15 ;
  wire \PCI-ROM/RB16 ;
  wire \PCI-ROM/RB17 ;
  wire \PCI-ROM/RB18 ;
  wire \PCI-ROM/RB19 ;
  wire \PCI-ROM/RB20 ;
  wire \PCI-ROM/RB21 ;
  wire \PCI-ROM/RB22 ;
  wire \PCI-ROM/RB23 ;
  wire \PCI-ROM/RB24 ;
  wire \PCI-ROM/RB25 ;
  wire \PCI-ROM/RB26 ;
  wire \PCI-ROM/RB27 ;
  wire \PCI-ROM/RB28 ;
  wire \PCI-ROM/RB29 ;
  wire \PCI-ROM/RB30 ;
  wire \PCI-ROM/RB31 ;
  wire \PCI-ROM/SEL2 ;
  wire \PCI-ROM/$1N8111 ;
  wire \PCI-ROM/SEL0 ;
  wire \PCI-ROM/$1N7806 ;
  wire \PCI-ROM/$1I7800/$1N2283 ;
  wire \PCI-ROM/$1I7800/$1N2277 ;
  wire \PCI-ROM/$1I7800/$1N2276 ;
  wire \PCI-ROM/$1I7800/$1N2275 ;
  wire \PCI-ROM/$1I8181/$1N2283 ;
  wire \PCI-ROM/$1I8181/$1N2277 ;
  wire \PCI-ROM/$1I8181/$1N2275 ;
  wire \PCI-ROM/$1I8225/$1N2277 ;
  wire \PCI-ROM/$1I8225/$1N2275 ;
  wire \PCI-ROM/$1I8276/$1N2277 ;
  wire \PCI-ROM/$1I8288/$1N2277 ;
  wire \PCI-ROM/$1I8332/$1N2290 ;
  wire \PCI-ROM/$1I8452/$1N2216 ;
  wire \$4I4029/$1N2778 ;
  wire \$4I4029/$1N2763 ;
  wire \$4I4029/ONE ;
  wire \$4I4029/EXP ;
  wire \$4I4029/$1N2759 ;
  wire \$4I4029/$1N2757 ;
  wire \$4I4029/$1N2755 ;
  wire \$4I4029/$1N2753 ;
  wire \$4I4029/$1N2751 ;
  wire \$4I4029/$1N2749 ;
  wire \$4I4029/$1N2734 ;
  wire \$4I4029/$1N2711 ;
  wire \$4I4029/$1N2616 ;
  wire \$4I4029/$1I2610/$1N86 ;
  wire \$4I4029/$1I2610/$1N87 ;
  wire \$4I4029/$1I2610/$1N81 ;
  wire \$4I4029/$1I2610/$1N82 ;
  wire \$4I4029/$1I2610/$1N71 ;
  wire \$4I4029/$1I2610/$1N70 ;
  wire \$4I4029/$1I2610/$1N66 ;
  wire \$4I4029/$1I2610/$1N65 ;
  wire \$4I4029/$1I2610/$1N61 ;
  wire \$4I4029/$1I2610/$1N62 ;
  wire \$4I4029/$1I2610/$1N56 ;
  wire \$4I4029/$1I2610/$1N55 ;
  wire \$4I4029/$1I2610/$1N51 ;
  wire \$4I4029/$1I2610/$1N50 ;
  wire \$4I4029/$1I2610/$1N48 ;
  wire \$4I4029/$1I2610/$1N45 ;
  wire \$4I4029/$1I2610/T7 ;
  wire \$4I4029/$1I2610/T3 ;
  wire \$4I4029/$1I2610/T2 ;
  wire \$4I4029/$1I2610/T5 ;
  wire \$4I4029/$1I2610/$1N20 ;
  wire \$4I4029/$1I2610/Q0 ;
  wire \$4I4029/$1I2610/Q1 ;
  wire \$4I4029/$1I2610/Q2 ;
  wire \$4I4029/$1I2610/Q3 ;
  wire \$4I4029/$1I2610/T6 ;
  wire \$4I4029/$1I2610/TC ;
  wire \$4I4029/$1I2610/T4 ;
  wire \$4I4029/$1I2610/Q4 ;
  wire \$4I4029/$1I2610/Q5 ;
  wire \$4I4029/$1I2610/Q6 ;
  wire \$4I4029/$1I2610/Q7 ;
  wire \$4I4029/$1I2610/$1I43/TQ ;
  wire \$4I4029/$1I2610/$1I43/MD ;
  wire \$4I4029/$1I2610/$1I43/$1I30/M1 ;
  wire \$4I4029/$1I2610/$1I43/$1I30/M0 ;
  wire \$4I4029/$1I2610/$1I44/$1N2216 ;
  wire \$4I4029/$1I2610/$1I47/$1N2216 ;
  wire \$4I4029/$1I2610/$1I49/$1N2216 ;
  wire \$4I4029/$1I2610/$1I52/$1N2216 ;
  wire \$4I4029/$1I2610/$1I53/TQ ;
  wire \$4I4029/$1I2610/$1I53/MD ;
  wire \$4I4029/$1I2610/$1I53/$1I30/M1 ;
  wire \$4I4029/$1I2610/$1I53/$1I30/M0 ;
  wire \$4I4029/$1I2610/$1I54/$1N2216 ;
  wire \$4I4029/$1I2610/$1I57/$1N2216 ;
  wire \$4I4029/$1I2610/$1I58/TQ ;
  wire \$4I4029/$1I2610/$1I58/MD ;
  wire \$4I4029/$1I2610/$1I58/$1I30/M1 ;
  wire \$4I4029/$1I2610/$1I58/$1I30/M0 ;
  wire \$4I4029/$1I2610/$1I59/TQ ;
  wire \$4I4029/$1I2610/$1I59/MD ;
  wire \$4I4029/$1I2610/$1I59/$1I30/M1 ;
  wire \$4I4029/$1I2610/$1I59/$1I30/M0 ;
  wire \$4I4029/$1I2610/$1I60/$1N2216 ;
  wire \$4I4029/$1I2610/$1I63/$1N2216 ;
  wire \$4I4029/$1I2610/$1I64/$1N2216 ;
  wire \$4I4029/$1I2610/$1I67/$1N2216 ;
  wire \$4I4029/$1I2610/$1I68/TQ ;
  wire \$4I4029/$1I2610/$1I68/MD ;
  wire \$4I4029/$1I2610/$1I68/$1I30/M1 ;
  wire \$4I4029/$1I2610/$1I68/$1I30/M0 ;
  wire \$4I4029/$1I2610/$1I69/$1N2216 ;
  wire \$4I4029/$1I2610/$1I72/$1N2216 ;
  wire \$4I4029/$1I2610/$1I73/TQ ;
  wire \$4I4029/$1I2610/$1I73/MD ;
  wire \$4I4029/$1I2610/$1I73/$1I30/M1 ;
  wire \$4I4029/$1I2610/$1I73/$1I30/M0 ;
  wire \$4I4029/$1I2610/$1I79/TQ ;
  wire \$4I4029/$1I2610/$1I79/MD ;
  wire \$4I4029/$1I2610/$1I79/$1I30/M1 ;
  wire \$4I4029/$1I2610/$1I79/$1I30/M0 ;
  wire \$4I4029/$1I2610/$1I80/$1N2216 ;
  wire \$4I4029/$1I2610/$1I83/$1N2216 ;
  wire \$4I4029/$1I2610/$1I84/TQ ;
  wire \$4I4029/$1I2610/$1I84/MD ;
  wire \$4I4029/$1I2610/$1I84/$1I30/M1 ;
  wire \$4I4029/$1I2610/$1I84/$1I30/M0 ;
  wire \$4I4029/$1I2610/$1I85/$1N2216 ;
  wire \$4I4029/$1I2610/$1I88/$1N2216 ;
  wire \$4I4029/$1I2615/$1N2216 ;
  wire \$4I4029/$1I2637/$1N86 ;
  wire \$4I4029/$1I2637/$1N87 ;
  wire \$4I4029/$1I2637/$1N81 ;
  wire \$4I4029/$1I2637/$1N82 ;
  wire \$4I4029/$1I2637/$1N71 ;
  wire \$4I4029/$1I2637/$1N70 ;
  wire \$4I4029/$1I2637/$1N66 ;
  wire \$4I4029/$1I2637/$1N65 ;
  wire \$4I4029/$1I2637/$1N61 ;
  wire \$4I4029/$1I2637/$1N62 ;
  wire \$4I4029/$1I2637/$1N56 ;
  wire \$4I4029/$1I2637/$1N55 ;
  wire \$4I4029/$1I2637/$1N51 ;
  wire \$4I4029/$1I2637/$1N50 ;
  wire \$4I4029/$1I2637/$1N48 ;
  wire \$4I4029/$1I2637/$1N45 ;
  wire \$4I4029/$1I2637/T7 ;
  wire \$4I4029/$1I2637/T3 ;
  wire \$4I4029/$1I2637/T2 ;
  wire \$4I4029/$1I2637/T5 ;
  wire \$4I4029/$1I2637/$1N20 ;
  wire \$4I4029/$1I2637/Q0 ;
  wire \$4I4029/$1I2637/Q1 ;
  wire \$4I4029/$1I2637/Q2 ;
  wire \$4I4029/$1I2637/Q3 ;
  wire \$4I4029/$1I2637/T6 ;
  wire \$4I4029/$1I2637/TC ;
  wire \$4I4029/$1I2637/T4 ;
  wire \$4I4029/$1I2637/Q4 ;
  wire \$4I4029/$1I2637/Q5 ;
  wire \$4I4029/$1I2637/Q6 ;
  wire \$4I4029/$1I2637/Q7 ;
  wire \$4I4029/$1I2637/$1I43/TQ ;
  wire \$4I4029/$1I2637/$1I43/MD ;
  wire \$4I4029/$1I2637/$1I43/$1I30/M1 ;
  wire \$4I4029/$1I2637/$1I43/$1I30/M0 ;
  wire \$4I4029/$1I2637/$1I44/$1N2216 ;
  wire \$4I4029/$1I2637/$1I47/$1N2216 ;
  wire \$4I4029/$1I2637/$1I49/$1N2216 ;
  wire \$4I4029/$1I2637/$1I52/$1N2216 ;
  wire \$4I4029/$1I2637/$1I53/TQ ;
  wire \$4I4029/$1I2637/$1I53/MD ;
  wire \$4I4029/$1I2637/$1I53/$1I30/M1 ;
  wire \$4I4029/$1I2637/$1I53/$1I30/M0 ;
  wire \$4I4029/$1I2637/$1I54/$1N2216 ;
  wire \$4I4029/$1I2637/$1I57/$1N2216 ;
  wire \$4I4029/$1I2637/$1I58/TQ ;
  wire \$4I4029/$1I2637/$1I58/MD ;
  wire \$4I4029/$1I2637/$1I58/$1I30/M1 ;
  wire \$4I4029/$1I2637/$1I58/$1I30/M0 ;
  wire \$4I4029/$1I2637/$1I59/TQ ;
  wire \$4I4029/$1I2637/$1I59/MD ;
  wire \$4I4029/$1I2637/$1I59/$1I30/M1 ;
  wire \$4I4029/$1I2637/$1I59/$1I30/M0 ;
  wire \$4I4029/$1I2637/$1I60/$1N2216 ;
  wire \$4I4029/$1I2637/$1I63/$1N2216 ;
  wire \$4I4029/$1I2637/$1I64/$1N2216 ;
  wire \$4I4029/$1I2637/$1I67/$1N2216 ;
  wire \$4I4029/$1I2637/$1I68/TQ ;
  wire \$4I4029/$1I2637/$1I68/MD ;
  wire \$4I4029/$1I2637/$1I68/$1I30/M1 ;
  wire \$4I4029/$1I2637/$1I68/$1I30/M0 ;
  wire \$4I4029/$1I2637/$1I69/$1N2216 ;
  wire \$4I4029/$1I2637/$1I72/$1N2216 ;
  wire \$4I4029/$1I2637/$1I73/TQ ;
  wire \$4I4029/$1I2637/$1I73/MD ;
  wire \$4I4029/$1I2637/$1I73/$1I30/M1 ;
  wire \$4I4029/$1I2637/$1I73/$1I30/M0 ;
  wire \$4I4029/$1I2637/$1I79/TQ ;
  wire \$4I4029/$1I2637/$1I79/MD ;
  wire \$4I4029/$1I2637/$1I79/$1I30/M1 ;
  wire \$4I4029/$1I2637/$1I79/$1I30/M0 ;
  wire \$4I4029/$1I2637/$1I80/$1N2216 ;
  wire \$4I4029/$1I2637/$1I83/$1N2216 ;
  wire \$4I4029/$1I2637/$1I84/TQ ;
  wire \$4I4029/$1I2637/$1I84/MD ;
  wire \$4I4029/$1I2637/$1I84/$1I30/M1 ;
  wire \$4I4029/$1I2637/$1I84/$1I30/M0 ;
  wire \$4I4029/$1I2637/$1I85/$1N2216 ;
  wire \$4I4029/$1I2637/$1I88/$1N2216 ;
  wire \$4I4029/$1I2645/$1N86 ;
  wire \$4I4029/$1I2645/$1N87 ;
  wire \$4I4029/$1I2645/$1N81 ;
  wire \$4I4029/$1I2645/$1N82 ;
  wire \$4I4029/$1I2645/$1N71 ;
  wire \$4I4029/$1I2645/$1N70 ;
  wire \$4I4029/$1I2645/$1N66 ;
  wire \$4I4029/$1I2645/$1N65 ;
  wire \$4I4029/$1I2645/$1N61 ;
  wire \$4I4029/$1I2645/$1N62 ;
  wire \$4I4029/$1I2645/$1N56 ;
  wire \$4I4029/$1I2645/$1N55 ;
  wire \$4I4029/$1I2645/$1N51 ;
  wire \$4I4029/$1I2645/$1N50 ;
  wire \$4I4029/$1I2645/$1N48 ;
  wire \$4I4029/$1I2645/$1N45 ;
  wire \$4I4029/$1I2645/T7 ;
  wire \$4I4029/$1I2645/T3 ;
  wire \$4I4029/$1I2645/T2 ;
  wire \$4I4029/$1I2645/T5 ;
  wire \$4I4029/$1I2645/$1N20 ;
  wire \$4I4029/$1I2645/Q0 ;
  wire \$4I4029/$1I2645/Q1 ;
  wire \$4I4029/$1I2645/Q2 ;
  wire \$4I4029/$1I2645/Q3 ;
  wire \$4I4029/$1I2645/T6 ;
  wire \$4I4029/$1I2645/TC ;
  wire \$4I4029/$1I2645/T4 ;
  wire \$4I4029/$1I2645/Q4 ;
  wire \$4I4029/$1I2645/Q5 ;
  wire \$4I4029/$1I2645/Q6 ;
  wire \$4I4029/$1I2645/Q7 ;
  wire \$4I4029/$1I2645/$1I43/TQ ;
  wire \$4I4029/$1I2645/$1I43/MD ;
  wire \$4I4029/$1I2645/$1I43/$1I30/M1 ;
  wire \$4I4029/$1I2645/$1I43/$1I30/M0 ;
  wire \$4I4029/$1I2645/$1I44/$1N2216 ;
  wire \$4I4029/$1I2645/$1I47/$1N2216 ;
  wire \$4I4029/$1I2645/$1I49/$1N2216 ;
  wire \$4I4029/$1I2645/$1I52/$1N2216 ;
  wire \$4I4029/$1I2645/$1I53/TQ ;
  wire \$4I4029/$1I2645/$1I53/MD ;
  wire \$4I4029/$1I2645/$1I53/$1I30/M1 ;
  wire \$4I4029/$1I2645/$1I53/$1I30/M0 ;
  wire \$4I4029/$1I2645/$1I54/$1N2216 ;
  wire \$4I4029/$1I2645/$1I57/$1N2216 ;
  wire \$4I4029/$1I2645/$1I58/TQ ;
  wire \$4I4029/$1I2645/$1I58/MD ;
  wire \$4I4029/$1I2645/$1I58/$1I30/M1 ;
  wire \$4I4029/$1I2645/$1I58/$1I30/M0 ;
  wire \$4I4029/$1I2645/$1I59/TQ ;
  wire \$4I4029/$1I2645/$1I59/MD ;
  wire \$4I4029/$1I2645/$1I59/$1I30/M1 ;
  wire \$4I4029/$1I2645/$1I59/$1I30/M0 ;
  wire \$4I4029/$1I2645/$1I60/$1N2216 ;
  wire \$4I4029/$1I2645/$1I63/$1N2216 ;
  wire \$4I4029/$1I2645/$1I64/$1N2216 ;
  wire \$4I4029/$1I2645/$1I67/$1N2216 ;
  wire \$4I4029/$1I2645/$1I68/TQ ;
  wire \$4I4029/$1I2645/$1I68/MD ;
  wire \$4I4029/$1I2645/$1I68/$1I30/M1 ;
  wire \$4I4029/$1I2645/$1I68/$1I30/M0 ;
  wire \$4I4029/$1I2645/$1I69/$1N2216 ;
  wire \$4I4029/$1I2645/$1I72/$1N2216 ;
  wire \$4I4029/$1I2645/$1I73/TQ ;
  wire \$4I4029/$1I2645/$1I73/MD ;
  wire \$4I4029/$1I2645/$1I73/$1I30/M1 ;
  wire \$4I4029/$1I2645/$1I73/$1I30/M0 ;
  wire \$4I4029/$1I2645/$1I79/TQ ;
  wire \$4I4029/$1I2645/$1I79/MD ;
  wire \$4I4029/$1I2645/$1I79/$1I30/M1 ;
  wire \$4I4029/$1I2645/$1I79/$1I30/M0 ;
  wire \$4I4029/$1I2645/$1I80/$1N2216 ;
  wire \$4I4029/$1I2645/$1I83/$1N2216 ;
  wire \$4I4029/$1I2645/$1I84/TQ ;
  wire \$4I4029/$1I2645/$1I84/MD ;
  wire \$4I4029/$1I2645/$1I84/$1I30/M1 ;
  wire \$4I4029/$1I2645/$1I84/$1I30/M0 ;
  wire \$4I4029/$1I2645/$1I85/$1N2216 ;
  wire \$4I4029/$1I2645/$1I88/$1N2216 ;
  wire \$4I4029/$1I2653/$1N86 ;
  wire \$4I4029/$1I2653/$1N87 ;
  wire \$4I4029/$1I2653/$1N81 ;
  wire \$4I4029/$1I2653/$1N82 ;
  wire \$4I4029/$1I2653/$1N71 ;
  wire \$4I4029/$1I2653/$1N70 ;
  wire \$4I4029/$1I2653/$1N66 ;
  wire \$4I4029/$1I2653/$1N65 ;
  wire \$4I4029/$1I2653/$1N61 ;
  wire \$4I4029/$1I2653/$1N62 ;
  wire \$4I4029/$1I2653/$1N56 ;
  wire \$4I4029/$1I2653/$1N55 ;
  wire \$4I4029/$1I2653/$1N51 ;
  wire \$4I4029/$1I2653/$1N50 ;
  wire \$4I4029/$1I2653/$1N48 ;
  wire \$4I4029/$1I2653/$1N45 ;
  wire \$4I4029/$1I2653/T7 ;
  wire \$4I4029/$1I2653/T3 ;
  wire \$4I4029/$1I2653/T2 ;
  wire \$4I4029/$1I2653/T5 ;
  wire \$4I4029/$1I2653/$1N20 ;
  wire \$4I4029/$1I2653/Q0 ;
  wire \$4I4029/$1I2653/Q1 ;
  wire \$4I4029/$1I2653/Q2 ;
  wire \$4I4029/$1I2653/Q3 ;
  wire \$4I4029/$1I2653/T6 ;
  wire \$4I4029/$1I2653/TC ;
  wire \$4I4029/$1I2653/T4 ;
  wire \$4I4029/$1I2653/Q4 ;
  wire \$4I4029/$1I2653/Q5 ;
  wire \$4I4029/$1I2653/Q6 ;
  wire \$4I4029/$1I2653/Q7 ;
  wire \$4I4029/$1I2653/$1I43/TQ ;
  wire \$4I4029/$1I2653/$1I43/MD ;
  wire \$4I4029/$1I2653/$1I43/$1I30/M1 ;
  wire \$4I4029/$1I2653/$1I43/$1I30/M0 ;
  wire \$4I4029/$1I2653/$1I44/$1N2216 ;
  wire \$4I4029/$1I2653/$1I47/$1N2216 ;
  wire \$4I4029/$1I2653/$1I49/$1N2216 ;
  wire \$4I4029/$1I2653/$1I52/$1N2216 ;
  wire \$4I4029/$1I2653/$1I53/TQ ;
  wire \$4I4029/$1I2653/$1I53/MD ;
  wire \$4I4029/$1I2653/$1I53/$1I30/M1 ;
  wire \$4I4029/$1I2653/$1I53/$1I30/M0 ;
  wire \$4I4029/$1I2653/$1I54/$1N2216 ;
  wire \$4I4029/$1I2653/$1I57/$1N2216 ;
  wire \$4I4029/$1I2653/$1I58/TQ ;
  wire \$4I4029/$1I2653/$1I58/MD ;
  wire \$4I4029/$1I2653/$1I58/$1I30/M1 ;
  wire \$4I4029/$1I2653/$1I58/$1I30/M0 ;
  wire \$4I4029/$1I2653/$1I59/TQ ;
  wire \$4I4029/$1I2653/$1I59/MD ;
  wire \$4I4029/$1I2653/$1I59/$1I30/M1 ;
  wire \$4I4029/$1I2653/$1I59/$1I30/M0 ;
  wire \$4I4029/$1I2653/$1I60/$1N2216 ;
  wire \$4I4029/$1I2653/$1I63/$1N2216 ;
  wire \$4I4029/$1I2653/$1I64/$1N2216 ;
  wire \$4I4029/$1I2653/$1I67/$1N2216 ;
  wire \$4I4029/$1I2653/$1I68/TQ ;
  wire \$4I4029/$1I2653/$1I68/MD ;
  wire \$4I4029/$1I2653/$1I68/$1I30/M1 ;
  wire \$4I4029/$1I2653/$1I68/$1I30/M0 ;
  wire \$4I4029/$1I2653/$1I69/$1N2216 ;
  wire \$4I4029/$1I2653/$1I72/$1N2216 ;
  wire \$4I4029/$1I2653/$1I73/TQ ;
  wire \$4I4029/$1I2653/$1I73/MD ;
  wire \$4I4029/$1I2653/$1I73/$1I30/M1 ;
  wire \$4I4029/$1I2653/$1I73/$1I30/M0 ;
  wire \$4I4029/$1I2653/$1I79/TQ ;
  wire \$4I4029/$1I2653/$1I79/MD ;
  wire \$4I4029/$1I2653/$1I79/$1I30/M1 ;
  wire \$4I4029/$1I2653/$1I79/$1I30/M0 ;
  wire \$4I4029/$1I2653/$1I80/$1N2216 ;
  wire \$4I4029/$1I2653/$1I83/$1N2216 ;
  wire \$4I4029/$1I2653/$1I84/TQ ;
  wire \$4I4029/$1I2653/$1I84/MD ;
  wire \$4I4029/$1I2653/$1I84/$1I30/M1 ;
  wire \$4I4029/$1I2653/$1I84/$1I30/M0 ;
  wire \$4I4029/$1I2653/$1I85/$1N2216 ;
  wire \$4I4029/$1I2653/$1I88/$1N2216 ;
  wire \$4I4029/$1I2661/$1N86 ;
  wire \$4I4029/$1I2661/$1N87 ;
  wire \$4I4029/$1I2661/$1N81 ;
  wire \$4I4029/$1I2661/$1N82 ;
  wire \$4I4029/$1I2661/$1N71 ;
  wire \$4I4029/$1I2661/$1N70 ;
  wire \$4I4029/$1I2661/$1N66 ;
  wire \$4I4029/$1I2661/$1N65 ;
  wire \$4I4029/$1I2661/$1N61 ;
  wire \$4I4029/$1I2661/$1N62 ;
  wire \$4I4029/$1I2661/$1N56 ;
  wire \$4I4029/$1I2661/$1N55 ;
  wire \$4I4029/$1I2661/$1N51 ;
  wire \$4I4029/$1I2661/$1N50 ;
  wire \$4I4029/$1I2661/$1N48 ;
  wire \$4I4029/$1I2661/$1N45 ;
  wire \$4I4029/$1I2661/T7 ;
  wire \$4I4029/$1I2661/T3 ;
  wire \$4I4029/$1I2661/T2 ;
  wire \$4I4029/$1I2661/T5 ;
  wire \$4I4029/$1I2661/$1N20 ;
  wire \$4I4029/$1I2661/Q0 ;
  wire \$4I4029/$1I2661/Q1 ;
  wire \$4I4029/$1I2661/Q2 ;
  wire \$4I4029/$1I2661/Q3 ;
  wire \$4I4029/$1I2661/T6 ;
  wire \$4I4029/$1I2661/TC ;
  wire \$4I4029/$1I2661/T4 ;
  wire \$4I4029/$1I2661/Q4 ;
  wire \$4I4029/$1I2661/Q5 ;
  wire \$4I4029/$1I2661/Q6 ;
  wire \$4I4029/$1I2661/Q7 ;
  wire \$4I4029/$1I2661/$1I43/TQ ;
  wire \$4I4029/$1I2661/$1I43/MD ;
  wire \$4I4029/$1I2661/$1I43/$1I30/M1 ;
  wire \$4I4029/$1I2661/$1I43/$1I30/M0 ;
  wire \$4I4029/$1I2661/$1I44/$1N2216 ;
  wire \$4I4029/$1I2661/$1I47/$1N2216 ;
  wire \$4I4029/$1I2661/$1I49/$1N2216 ;
  wire \$4I4029/$1I2661/$1I52/$1N2216 ;
  wire \$4I4029/$1I2661/$1I53/TQ ;
  wire \$4I4029/$1I2661/$1I53/MD ;
  wire \$4I4029/$1I2661/$1I53/$1I30/M1 ;
  wire \$4I4029/$1I2661/$1I53/$1I30/M0 ;
  wire \$4I4029/$1I2661/$1I54/$1N2216 ;
  wire \$4I4029/$1I2661/$1I57/$1N2216 ;
  wire \$4I4029/$1I2661/$1I58/TQ ;
  wire \$4I4029/$1I2661/$1I58/MD ;
  wire \$4I4029/$1I2661/$1I58/$1I30/M1 ;
  wire \$4I4029/$1I2661/$1I58/$1I30/M0 ;
  wire \$4I4029/$1I2661/$1I59/TQ ;
  wire \$4I4029/$1I2661/$1I59/MD ;
  wire \$4I4029/$1I2661/$1I59/$1I30/M1 ;
  wire \$4I4029/$1I2661/$1I59/$1I30/M0 ;
  wire \$4I4029/$1I2661/$1I60/$1N2216 ;
  wire \$4I4029/$1I2661/$1I63/$1N2216 ;
  wire \$4I4029/$1I2661/$1I64/$1N2216 ;
  wire \$4I4029/$1I2661/$1I67/$1N2216 ;
  wire \$4I4029/$1I2661/$1I68/TQ ;
  wire \$4I4029/$1I2661/$1I68/MD ;
  wire \$4I4029/$1I2661/$1I68/$1I30/M1 ;
  wire \$4I4029/$1I2661/$1I68/$1I30/M0 ;
  wire \$4I4029/$1I2661/$1I69/$1N2216 ;
  wire \$4I4029/$1I2661/$1I72/$1N2216 ;
  wire \$4I4029/$1I2661/$1I73/TQ ;
  wire \$4I4029/$1I2661/$1I73/MD ;
  wire \$4I4029/$1I2661/$1I73/$1I30/M1 ;
  wire \$4I4029/$1I2661/$1I73/$1I30/M0 ;
  wire \$4I4029/$1I2661/$1I79/TQ ;
  wire \$4I4029/$1I2661/$1I79/MD ;
  wire \$4I4029/$1I2661/$1I79/$1I30/M1 ;
  wire \$4I4029/$1I2661/$1I79/$1I30/M0 ;
  wire \$4I4029/$1I2661/$1I80/$1N2216 ;
  wire \$4I4029/$1I2661/$1I83/$1N2216 ;
  wire \$4I4029/$1I2661/$1I84/TQ ;
  wire \$4I4029/$1I2661/$1I84/MD ;
  wire \$4I4029/$1I2661/$1I84/$1I30/M1 ;
  wire \$4I4029/$1I2661/$1I84/$1I30/M0 ;
  wire \$4I4029/$1I2661/$1I85/$1N2216 ;
  wire \$4I4029/$1I2661/$1I88/$1N2216 ;
  wire \$4I4029/$1I2730/$1N2216 ;
  wire \$4I4076/$1N2216 ;
  wire \$4I4095/$1N2216 ;
  wire \$4I4096/$1N2216 ;
  wire \$4I4097/$1N2216 ;
  wire \$4I4098/$1N2216 ;
  wire \$4I4099/$1N2216 ;
  wire \$4I4100/$1N2216 ;
  wire \$4I4101/$1N2216 ;
  wire \$4I4102/$1N2216 ;
  wire \$4I4103/$1N2216 ;
  wire \OEADI/$1N4030 ;
  wire \OEADI/$1N4036 ;
  wire \OEADI/$1N4042 ;
  wire \OEADI/OAI64_0 ;
  wire \OEADI/OAI64_1 ;
  wire \OEADI/MIDDLE ;
  wire \OEADI/$1N3986 ;
  wire \OEADI/OAI32_1 ;
  wire \OEADI/OAI32_0 ;
  wire \OEADI/CFG_SELFQ ;
  wire \OEADI/$1N3857 ;
  wire \OEADI/$1N3855 ;
  wire \OEADI/M_DATAQ ;
  wire \$5I3771/M1 ;
  wire \$5I3771/M0 ;
  wire \$5I3778/$1N2216 ;
  wire \$5I3781/M1 ;
  wire \$5I3781/M0 ;
  wire \$5I3782/$1N2216 ;
  wire \DEVSEL/$1N2307 ;
  wire \DEVSEL/D1_9541 ;
  wire \DEVSEL/D3_9540 ;
  wire \DEVSEL/D2_9539 ;
  wire \DEVSEL/IN ;
  wire \DEVSEL/$1N2275 ;
  wire \DEVSEL/$1I2276/$1N2216 ;
  wire \DEVSEL/$1I2306/$1N2216 ;
  wire \DEVSEL/$1I2310/M23 ;
  wire \DEVSEL/$1I2310/M01 ;
  wire \DEVSEL/$1I2310/M01/M0 ;
  wire \DEVSEL/$1I2310/M01/M1 ;
  wire \DEVSEL/$1I2310/M23/M0 ;
  wire \DEVSEL/$1I2310/M23/M1 ;
  wire \ACK64/$1N2307 ;
  wire \ACK64/D1_9585 ;
  wire \ACK64/D3_9584 ;
  wire \ACK64/D2_9583 ;
  wire \ACK64/IN ;
  wire \ACK64/$1N2275 ;
  wire \ACK64/$1I2276/$1N2216 ;
  wire \ACK64/$1I2306/$1N2216 ;
  wire \ACK64/$1I2310/M23 ;
  wire \ACK64/$1I2310/M01 ;
  wire \ACK64/$1I2310/M01/M0 ;
  wire \ACK64/$1I2310/M01/M1 ;
  wire \ACK64/$1I2310/M23/M0 ;
  wire \ACK64/$1I2310/M23/M1 ;
  wire \FRAME/$1N2307 ;
  wire \FRAME/D1_9629 ;
  wire \FRAME/D3_9628 ;
  wire \FRAME/D2_9627 ;
  wire \FRAME/IN ;
  wire \FRAME/$1N2275 ;
  wire \FRAME/$1I2276/$1N2216 ;
  wire \FRAME/$1I2306/$1N2216 ;
  wire \FRAME/$1I2310/M23 ;
  wire \FRAME/$1I2310/M01 ;
  wire \FRAME/$1I2310/M01/M0 ;
  wire \FRAME/$1I2310/M01/M1 ;
  wire \FRAME/$1I2310/M23/M0 ;
  wire \FRAME/$1I2310/M23/M1 ;
  wire \$6I1174/$1N2216 ;
  wire \TRDY/$1N2307 ;
  wire \TRDY/D1_9675 ;
  wire \TRDY/D3_9674 ;
  wire \TRDY/D2_9673 ;
  wire \TRDY/IN ;
  wire \TRDY/$1N2275 ;
  wire \TRDY/$1I2276/$1N2216 ;
  wire \TRDY/$1I2306/$1N2216 ;
  wire \TRDY/$1I2310/M23 ;
  wire \TRDY/$1I2310/M01 ;
  wire \TRDY/$1I2310/M01/M0 ;
  wire \TRDY/$1I2310/M01/M1 ;
  wire \TRDY/$1I2310/M23/M0 ;
  wire \TRDY/$1I2310/M23/M1 ;
  wire \REQ64/$1N2307 ;
  wire \REQ64/D1_9719 ;
  wire \REQ64/D3_9718 ;
  wire \REQ64/D2_9717 ;
  wire \REQ64/IN ;
  wire \REQ64/$1N2275 ;
  wire \REQ64/$1I2276/$1N2216 ;
  wire \REQ64/$1I2306/$1N2216 ;
  wire \REQ64/$1I2310/M23 ;
  wire \REQ64/$1I2310/M01 ;
  wire \REQ64/$1I2310/M01/M0 ;
  wire \REQ64/$1I2310/M01/M1 ;
  wire \REQ64/$1I2310/M23/M0 ;
  wire \REQ64/$1I2310/M23/M1 ;
  wire \IRDY/$1N2307 ;
  wire \IRDY/D1_9763 ;
  wire \IRDY/D3_9762 ;
  wire \IRDY/D2_9761 ;
  wire \IRDY/IN ;
  wire \IRDY/$1N2275 ;
  wire \IRDY/$1I2276/$1N2216 ;
  wire \IRDY/$1I2306/$1N2216 ;
  wire \IRDY/$1I2310/M23 ;
  wire \IRDY/$1I2310/M01 ;
  wire \IRDY/$1I2310/M01/M0 ;
  wire \IRDY/$1I2310/M01/M1 ;
  wire \IRDY/$1I2310/M23/M0 ;
  wire \IRDY/$1I2310/M23/M1 ;
  wire \STOP/$1N2307 ;
  wire \STOP/D1_9807 ;
  wire \STOP/D3_9806 ;
  wire \STOP/D2_9805 ;
  wire \STOP/IN ;
  wire \STOP/$1N2275 ;
  wire \STOP/$1I2276/$1N2216 ;
  wire \STOP/$1I2306/$1N2216 ;
  wire \STOP/$1I2310/M23 ;
  wire \STOP/$1I2310/M01 ;
  wire \STOP/$1I2310/M01/M0 ;
  wire \STOP/$1I2310/M01/M1 ;
  wire \STOP/$1I2310/M23/M0 ;
  wire \STOP/$1I2310/M23/M1 ;
  wire \PERR/$1N2286 ;
  wire \PERR/$1N2289 ;
  wire \PERR/$1I2285/$1N2216 ;
  wire \PERR/$1I2288/$1N2216 ;
  wire \SERR/$1N2286 ;
  wire \SERR/$1N2289 ;
  wire \SERR/$1I2285/$1N2216 ;
  wire \SERR/$1I2288/$1N2216 ;
  wire \$6I950/$1N2216 ;
  wire \IDSEL/$1N2286 ;
  wire \IDSEL/$1N2289 ;
  wire \IDSEL/$1I2285/$1N2216 ;
  wire \IDSEL/$1I2288/$1N2216 ;
  wire \$6I961/$1N2216 ;
  wire \$7I576/M1 ;
  wire \$7I576/M0 ;
  wire \$7I577/M1 ;
  wire \$7I577/M0 ;
  wire \$7I580/$1N2283 ;
  wire \$7I580/$1N2277 ;
  wire \$7I580/$1N2276 ;
  wire \$7I580/$1N2275 ;
  wire \$7I622/M1 ;
  wire \$7I622/M0 ;
  wire \$7I623/M1 ;
  wire \$7I623/M0 ;
  wire \$7I632/$1N2216 ;
  wire \$7I633/$1N2216 ;
  wire \$7I746/$1N2216 ;
  wire \$7I824/M1 ;
  wire \$7I824/M0 ;
  wire \$7I826/M1 ;
  wire \$7I826/M0 ;
  wire \$7I828/M1 ;
  wire \$7I828/M0 ;
  wire \$7I830/M1 ;
  wire \$7I830/M0 ;
  wire \$7I832/M1 ;
  wire \$7I832/M0 ;
  wire \$7I834/M1 ;
  wire \$7I834/M0 ;
  wire \$7I836/M1 ;
  wire \$7I836/M0 ;
  wire \$7I838/M1 ;
  wire \$7I838/M0 ;
  wire \$7I861/$1N2216 ;
  wire \$7I862/$1N2216 ;
  wire \PCI-CBE/$1N2786 ;
  wire \PCI-CBE/SWITCH ;
  wire \PCI-CBE/TO_SW ;
  wire \PCI-CBE/TO_ACK ;
  wire \PCI-CBE/IO3/$1N2321 ;
  wire \PCI-CBE/IO3/D_SLO ;
  wire \PCI-CBE/IO3/$1I2296/M1 ;
  wire \PCI-CBE/IO3/$1I2296/M0 ;
  wire \PCI-CBE/IO3/$1I2303/M1 ;
  wire \PCI-CBE/IO3/$1I2303/M0 ;
  wire \PCI-CBE/IO2/$1N2321 ;
  wire \PCI-CBE/IO2/D_SLO ;
  wire \PCI-CBE/IO2/$1I2296/M1 ;
  wire \PCI-CBE/IO2/$1I2296/M0 ;
  wire \PCI-CBE/IO2/$1I2303/M1 ;
  wire \PCI-CBE/IO2/$1I2303/M0 ;
  wire \PCI-CBE/IO1/$1N2321 ;
  wire \PCI-CBE/IO1/D_SLO ;
  wire \PCI-CBE/IO1/$1I2296/M1 ;
  wire \PCI-CBE/IO1/$1I2296/M0 ;
  wire \PCI-CBE/IO1/$1I2303/M1 ;
  wire \PCI-CBE/IO1/$1I2303/M0 ;
  wire \PCI-CBE/IO0/$1N2321 ;
  wire \PCI-CBE/IO0/D_SLO ;
  wire \PCI-CBE/IO0/$1I2296/M1 ;
  wire \PCI-CBE/IO0/$1I2296/M0 ;
  wire \PCI-CBE/IO0/$1I2303/M1 ;
  wire \PCI-CBE/IO0/$1I2303/M0 ;
  wire \PCI-CBE/$1I2777/M1 ;
  wire \PCI-CBE/$1I2777/M0 ;
  wire \PCI-CBE/$1I2779/M1 ;
  wire \PCI-CBE/$1I2779/M0 ;
  wire \PCI-CBE/$1I2787/$1N2216 ;
  wire \PCI-AD/D_SLO0 ;
  wire \PCI-AD/D_SLO1 ;
  wire \PCI-AD/D_SLO2 ;
  wire \PCI-AD/D_SLO3 ;
  wire \PCI-AD/D_SLO8 ;
  wire \PCI-AD/D_SLO9 ;
  wire \PCI-AD/D_SLO10 ;
  wire \PCI-AD/D_SLO11 ;
  wire \PCI-AD/D_SLO16 ;
  wire \PCI-AD/D_SLO17 ;
  wire \PCI-AD/D_SLO18 ;
  wire \PCI-AD/D_SLO19 ;
  wire \PCI-AD/D_SLO24 ;
  wire \PCI-AD/D_SLO25 ;
  wire \PCI-AD/D_SLO26 ;
  wire \PCI-AD/D_SLO27 ;
  wire \PCI-AD/D_SLO7 ;
  wire \PCI-AD/D_SLO5 ;
  wire \PCI-AD/D_SLO6 ;
  wire \PCI-AD/D_SLO4 ;
  wire \PCI-AD/D_SLO15 ;
  wire \PCI-AD/D_SLO13 ;
  wire \PCI-AD/D_SLO14 ;
  wire \PCI-AD/D_SLO12 ;
  wire \PCI-AD/D_SLO23 ;
  wire \PCI-AD/D_SLO21 ;
  wire \PCI-AD/D_SLO22 ;
  wire \PCI-AD/D_SLO20 ;
  wire \PCI-AD/D_SLO31 ;
  wire \PCI-AD/D_SLO29 ;
  wire \PCI-AD/D_SLO30 ;
  wire \PCI-AD/D_SLO28 ;
  wire \PCI-AD/IO28/$1I2246/M1 ;
  wire \PCI-AD/IO28/$1I2246/M0 ;
  wire \PCI-AD/IO30/$1I2246/M1 ;
  wire \PCI-AD/IO30/$1I2246/M0 ;
  wire \PCI-AD/IO29/$1I2246/M1 ;
  wire \PCI-AD/IO29/$1I2246/M0 ;
  wire \PCI-AD/IO31/$1I2246/M1 ;
  wire \PCI-AD/IO31/$1I2246/M0 ;
  wire \PCI-AD/IO20/$1I2246/M1 ;
  wire \PCI-AD/IO20/$1I2246/M0 ;
  wire \PCI-AD/IO22/$1I2246/M1 ;
  wire \PCI-AD/IO22/$1I2246/M0 ;
  wire \PCI-AD/IO21/$1I2246/M1 ;
  wire \PCI-AD/IO21/$1I2246/M0 ;
  wire \PCI-AD/IO23/$1I2246/M1 ;
  wire \PCI-AD/IO23/$1I2246/M0 ;
  wire \PCI-AD/IO12/$1I2246/M1 ;
  wire \PCI-AD/IO12/$1I2246/M0 ;
  wire \PCI-AD/IO14/$1I2246/M1 ;
  wire \PCI-AD/IO14/$1I2246/M0 ;
  wire \PCI-AD/IO13/$1I2246/M1 ;
  wire \PCI-AD/IO13/$1I2246/M0 ;
  wire \PCI-AD/IO15/$1I2246/M1 ;
  wire \PCI-AD/IO15/$1I2246/M0 ;
  wire \PCI-AD/IO4/$1I2246/M1 ;
  wire \PCI-AD/IO4/$1I2246/M0 ;
  wire \PCI-AD/IO6/$1I2246/M1 ;
  wire \PCI-AD/IO6/$1I2246/M0 ;
  wire \PCI-AD/IO5/$1I2246/M1 ;
  wire \PCI-AD/IO5/$1I2246/M0 ;
  wire \PCI-AD/IO7/$1I2246/M1 ;
  wire \PCI-AD/IO7/$1I2246/M0 ;
  wire \PCI-AD/$1I2927/M1 ;
  wire \PCI-AD/$1I2927/M0 ;
  wire \PCI-AD/$1I2928/M1 ;
  wire \PCI-AD/$1I2928/M0 ;
  wire \PCI-AD/$1I2929/M1 ;
  wire \PCI-AD/$1I2929/M0 ;
  wire \PCI-AD/$1I2930/M1 ;
  wire \PCI-AD/$1I2930/M0 ;
  wire \PCI-AD/$1I2931/M1 ;
  wire \PCI-AD/$1I2931/M0 ;
  wire \PCI-AD/$1I2932/M1 ;
  wire \PCI-AD/$1I2932/M0 ;
  wire \PCI-AD/$1I2933/M1 ;
  wire \PCI-AD/$1I2933/M0 ;
  wire \PCI-AD/$1I2934/M1 ;
  wire \PCI-AD/$1I2934/M0 ;
  wire \PCI-AD/$1I2935/M1 ;
  wire \PCI-AD/$1I2935/M0 ;
  wire \PCI-AD/$1I2936/M1 ;
  wire \PCI-AD/$1I2936/M0 ;
  wire \PCI-AD/$1I2937/M1 ;
  wire \PCI-AD/$1I2937/M0 ;
  wire \PCI-AD/$1I2938/M1 ;
  wire \PCI-AD/$1I2938/M0 ;
  wire \PCI-AD/$1I2939/M1 ;
  wire \PCI-AD/$1I2939/M0 ;
  wire \PCI-AD/$1I2940/M1 ;
  wire \PCI-AD/$1I2940/M0 ;
  wire \PCI-AD/$1I2941/M1 ;
  wire \PCI-AD/$1I2941/M0 ;
  wire \PCI-AD/$1I2942/M1 ;
  wire \PCI-AD/$1I2942/M0 ;
  wire \PCI-AD/$1I2943/M1 ;
  wire \PCI-AD/$1I2943/M0 ;
  wire \PCI-AD/$1I2944/M1 ;
  wire \PCI-AD/$1I2944/M0 ;
  wire \PCI-AD/$1I2945/M1 ;
  wire \PCI-AD/$1I2945/M0 ;
  wire \PCI-AD/$1I2946/M1 ;
  wire \PCI-AD/$1I2946/M0 ;
  wire \PCI-AD/$1I2947/M1 ;
  wire \PCI-AD/$1I2947/M0 ;
  wire \PCI-AD/$1I2948/M1 ;
  wire \PCI-AD/$1I2948/M0 ;
  wire \PCI-AD/$1I2949/M1 ;
  wire \PCI-AD/$1I2949/M0 ;
  wire \PCI-AD/$1I2950/M1 ;
  wire \PCI-AD/$1I2950/M0 ;
  wire \PCI-AD/$1I2951/M1 ;
  wire \PCI-AD/$1I2951/M0 ;
  wire \PCI-AD/$1I2952/M1 ;
  wire \PCI-AD/$1I2952/M0 ;
  wire \PCI-AD/$1I2953/M1 ;
  wire \PCI-AD/$1I2953/M0 ;
  wire \PCI-AD/$1I2954/M1 ;
  wire \PCI-AD/$1I2954/M0 ;
  wire \PCI-AD/$1I2955/M1 ;
  wire \PCI-AD/$1I2955/M0 ;
  wire \PCI-AD/$1I2956/M1 ;
  wire \PCI-AD/$1I2956/M0 ;
  wire \PCI-AD/$1I2957/M1 ;
  wire \PCI-AD/$1I2957/M0 ;
  wire \PCI-AD/$1I2958/M1 ;
  wire \PCI-AD/$1I2958/M0 ;
  wire \PCI-AD/IO27/$1I2246/M1 ;
  wire \PCI-AD/IO27/$1I2246/M0 ;
  wire \PCI-AD/IO26/$1I2246/M1 ;
  wire \PCI-AD/IO26/$1I2246/M0 ;
  wire \PCI-AD/IO25/$1I2246/M1 ;
  wire \PCI-AD/IO25/$1I2246/M0 ;
  wire \PCI-AD/IO24/$1I2246/M1 ;
  wire \PCI-AD/IO24/$1I2246/M0 ;
  wire \PCI-AD/IO19/$1I2246/M1 ;
  wire \PCI-AD/IO19/$1I2246/M0 ;
  wire \PCI-AD/IO18/$1I2246/M1 ;
  wire \PCI-AD/IO18/$1I2246/M0 ;
  wire \PCI-AD/IO17/$1I2246/M1 ;
  wire \PCI-AD/IO17/$1I2246/M0 ;
  wire \PCI-AD/IO16/$1I2246/M1 ;
  wire \PCI-AD/IO16/$1I2246/M0 ;
  wire \PCI-AD/IO11/$1I2246/M1 ;
  wire \PCI-AD/IO11/$1I2246/M0 ;
  wire \PCI-AD/IO10/$1I2246/M1 ;
  wire \PCI-AD/IO10/$1I2246/M0 ;
  wire \PCI-AD/IO9/$1I2246/M1 ;
  wire \PCI-AD/IO9/$1I2246/M0 ;
  wire \PCI-AD/IO8/$1I2246/M1 ;
  wire \PCI-AD/IO8/$1I2246/M0 ;
  wire \PCI-AD/IO3/$1I2246/M1 ;
  wire \PCI-AD/IO3/$1I2246/M0 ;
  wire \PCI-AD/IO2/$1I2246/M1 ;
  wire \PCI-AD/IO2/$1I2246/M0 ;
  wire \PCI-AD/IO1/$1I2246/M1 ;
  wire \PCI-AD/IO1/$1I2246/M0 ;
  wire \PCI-AD/IO0/$1I2246/M1 ;
  wire \PCI-AD/IO0/$1I2246/M0 ;
  wire \PCI-AD64/IO28/$1I2246/M1 ;
  wire \PCI-AD64/IO28/$1I2246/M0 ;
  wire \PCI-AD64/IO30/$1I2246/M1 ;
  wire \PCI-AD64/IO30/$1I2246/M0 ;
  wire \PCI-AD64/IO29/$1I2246/M1 ;
  wire \PCI-AD64/IO29/$1I2246/M0 ;
  wire \PCI-AD64/IO31/$1I2246/M1 ;
  wire \PCI-AD64/IO31/$1I2246/M0 ;
  wire \PCI-AD64/IO20/$1I2246/M1 ;
  wire \PCI-AD64/IO20/$1I2246/M0 ;
  wire \PCI-AD64/IO22/$1I2246/M1 ;
  wire \PCI-AD64/IO22/$1I2246/M0 ;
  wire \PCI-AD64/IO21/$1I2246/M1 ;
  wire \PCI-AD64/IO21/$1I2246/M0 ;
  wire \PCI-AD64/IO23/$1I2246/M1 ;
  wire \PCI-AD64/IO23/$1I2246/M0 ;
  wire \PCI-AD64/IO12/$1I2246/M1 ;
  wire \PCI-AD64/IO12/$1I2246/M0 ;
  wire \PCI-AD64/IO14/$1I2246/M1 ;
  wire \PCI-AD64/IO14/$1I2246/M0 ;
  wire \PCI-AD64/IO13/$1I2246/M1 ;
  wire \PCI-AD64/IO13/$1I2246/M0 ;
  wire \PCI-AD64/IO15/$1I2246/M1 ;
  wire \PCI-AD64/IO15/$1I2246/M0 ;
  wire \PCI-AD64/IO4/$1I2246/M1 ;
  wire \PCI-AD64/IO4/$1I2246/M0 ;
  wire \PCI-AD64/IO6/$1I2246/M1 ;
  wire \PCI-AD64/IO6/$1I2246/M0 ;
  wire \PCI-AD64/IO5/$1I2246/M1 ;
  wire \PCI-AD64/IO5/$1I2246/M0 ;
  wire \PCI-AD64/IO7/$1I2246/M1 ;
  wire \PCI-AD64/IO7/$1I2246/M0 ;
  wire \PCI-AD64/IO27/$1I2246/M1 ;
  wire \PCI-AD64/IO27/$1I2246/M0 ;
  wire \PCI-AD64/IO26/$1I2246/M1 ;
  wire \PCI-AD64/IO26/$1I2246/M0 ;
  wire \PCI-AD64/IO25/$1I2246/M1 ;
  wire \PCI-AD64/IO25/$1I2246/M0 ;
  wire \PCI-AD64/IO24/$1I2246/M1 ;
  wire \PCI-AD64/IO24/$1I2246/M0 ;
  wire \PCI-AD64/IO19/$1I2246/M1 ;
  wire \PCI-AD64/IO19/$1I2246/M0 ;
  wire \PCI-AD64/IO18/$1I2246/M1 ;
  wire \PCI-AD64/IO18/$1I2246/M0 ;
  wire \PCI-AD64/IO17/$1I2246/M1 ;
  wire \PCI-AD64/IO17/$1I2246/M0 ;
  wire \PCI-AD64/IO16/$1I2246/M1 ;
  wire \PCI-AD64/IO16/$1I2246/M0 ;
  wire \PCI-AD64/IO11/$1I2246/M1 ;
  wire \PCI-AD64/IO11/$1I2246/M0 ;
  wire \PCI-AD64/IO10/$1I2246/M1 ;
  wire \PCI-AD64/IO10/$1I2246/M0 ;
  wire \PCI-AD64/IO9/$1I2246/M1 ;
  wire \PCI-AD64/IO9/$1I2246/M0 ;
  wire \PCI-AD64/IO8/$1I2246/M1 ;
  wire \PCI-AD64/IO8/$1I2246/M0 ;
  wire \PCI-AD64/IO3/$1I2246/M1 ;
  wire \PCI-AD64/IO3/$1I2246/M0 ;
  wire \PCI-AD64/IO2/$1I2246/M1 ;
  wire \PCI-AD64/IO2/$1I2246/M0 ;
  wire \PCI-AD64/IO1/$1I2246/M1 ;
  wire \PCI-AD64/IO1/$1I2246/M0 ;
  wire \PCI-AD64/IO0/$1I2246/M1 ;
  wire \PCI-AD64/IO0/$1I2246/M0 ;
  wire \PCI-CBE64/$1N2781 ;
  wire \PCI-CBE64/$1N2783 ;
  wire \PCI-CBE64/$1N2779 ;
  wire \PCI-CBE64/$1N2787 ;
  wire \PCI-CBE64/$1N2789 ;
  wire \PCI-CBE64/$1N2785 ;
  wire \PCI-CBE64/$1N2793 ;
  wire \PCI-CBE64/$1N2795 ;
  wire \PCI-CBE64/$1N2791 ;
  wire \PCI-CBE64/$1N2799 ;
  wire \PCI-CBE64/$1N2801 ;
  wire \PCI-CBE64/$1N2797 ;
  wire \PCI-CBE64/IO3/$1N2321 ;
  wire \PCI-CBE64/IO3/D_SLO ;
  wire \PCI-CBE64/IO3/$1I2296/M1 ;
  wire \PCI-CBE64/IO3/$1I2296/M0 ;
  wire \PCI-CBE64/IO3/$1I2303/M1 ;
  wire \PCI-CBE64/IO3/$1I2303/M0 ;
  wire \PCI-CBE64/IO2/$1N2321 ;
  wire \PCI-CBE64/IO2/D_SLO ;
  wire \PCI-CBE64/IO2/$1I2296/M1 ;
  wire \PCI-CBE64/IO2/$1I2296/M0 ;
  wire \PCI-CBE64/IO2/$1I2303/M1 ;
  wire \PCI-CBE64/IO2/$1I2303/M0 ;
  wire \PCI-CBE64/IO1/$1N2321 ;
  wire \PCI-CBE64/IO1/D_SLO ;
  wire \PCI-CBE64/IO1/$1I2296/M1 ;
  wire \PCI-CBE64/IO1/$1I2296/M0 ;
  wire \PCI-CBE64/IO1/$1I2303/M1 ;
  wire \PCI-CBE64/IO1/$1I2303/M0 ;
  wire \PCI-CBE64/IO0/$1N2321 ;
  wire \PCI-CBE64/IO0/D_SLO ;
  wire \PCI-CBE64/IO0/$1I2296/M1 ;
  wire \PCI-CBE64/IO0/$1I2296/M0 ;
  wire \PCI-CBE64/IO0/$1I2303/M1 ;
  wire \PCI-CBE64/IO0/$1I2303/M0 ;
  wire \PCI-CBE64/$1I2777/$1N2216 ;
  wire \PCI-CBE64/$1I2780/$1N2216 ;
  wire \PCI-CBE64/$1I2782/$1N2216 ;
  wire \PCI-CBE64/$1I2784/$1N2216 ;
  wire \PCI-CBE64/$1I2786/$1N2216 ;
  wire \PCI-CBE64/$1I2788/$1N2216 ;
  wire \PCI-CBE64/$1I2790/$1N2216 ;
  wire \PCI-CBE64/$1I2792/$1N2216 ;
  wire \PCI-CBE64/$1I2794/$1N2216 ;
  wire \PCI-CBE64/$1I2796/$1N2216 ;
  wire \PCI-CBE64/$1I2798/$1N2216 ;
  wire \PCI-CBE64/$1I2800/$1N2216 ;
  wire \NlwInverterSignal_$3I3487/I0 ;
  wire \NlwInverterSignal_$3I3492/I0 ;
  wire \NlwInverterSignal_$3I3496/I0 ;
  wire \NlwInverterSignal_$4I4017/I0 ;
  wire \NlwInverterSignal_$4I4017/I1 ;
  wire \NlwInverterSignal_$4I4017/O ;
  wire \NlwInverterSignal_$6I1168/I0 ;
  wire \NlwInverterSignal_$6I1168/I1 ;
  wire \NlwInverterSignal_$6I1169/I0 ;
  wire \NlwInverterSignal_$6I1170/I0 ;
  wire \NlwInverterSignal_$6I1172/I0 ;
  wire \NlwInverterSignal_$7I129/I0 ;
  wire \NlwInverterSignal_$7I129/I1 ;
  wire \NlwInverterSignal_$7I130/I0 ;
  wire \NlwInverterSignal_$7I131/I0 ;
  wire \NlwInverterSignal_$7I132/I0 ;
  wire \NlwInverterSignal_$7I132/I1 ;
  wire \NlwInverterSignal_$7I133/I0 ;
  wire \NlwInverterSignal_$7I133/I1 ;
  wire \NlwInverterSignal_$7I133/I2 ;
  wire \NlwInverterSignal_$7I134/I0 ;
  wire \NlwInverterSignal_$7I141/I0 ;
  wire \NlwInverterSignal_$7I141/I1 ;
  wire VCC;
  wire GND;
  wire \NlwInverterSignal_$7I863/I0 ;
  wire \NlwInverterSignal_MASTER/$4I3271/I0 ;
  wire \NlwInverterSignal_MASTER/$4I3271/I1 ;
  wire \NlwInverterSignal_MASTER/$4I3271/I2 ;
  wire \NlwInverterSignal_MASTER/$4I3102/I0 ;
  wire \NlwInverterSignal_MASTER/$4I3102/I1 ;
  wire \NlwInverterSignal_MASTER/$4I3072/I0 ;
  wire \NlwInverterSignal_MASTER/$4I3051/I0 ;
  wire \NlwInverterSignal_MASTER/$4I2686/I0 ;
  wire \NlwInverterSignal_MASTER/$4I2686/I1 ;
  wire \NlwInverterSignal_MASTER/$4I2686/I2 ;
  wire \NlwInverterSignal_MASTER/I_IDLE/$1I2807/I0 ;
  wire \NlwInverterSignal_MASTER/I_IDLE/$1I2715/I0 ;
  wire \NlwInverterSignal_MASTER/I_IDLE/$1I2715/I1 ;
  wire \NlwInverterSignal_MASTER/I_IDLE/$1I2715/O ;
  wire \NlwInverterSignal_MASTER/I_IDLE/$1I2647/I0 ;
  wire \NlwInverterSignal_MASTER/I_IDLE/$1I2594/I0 ;
  wire \NlwInverterSignal_MASTER/I_IDLE/$1I2593/I0 ;
  wire \NlwInverterSignal_MASTER/ADDR/$1I2632/I0 ;
  wire \NlwInverterSignal_MASTER/ADDR/$1I2630/O ;
  wire \NlwInverterSignal_MASTER/ADDR/$1I2623/I0 ;
  wire \NlwInverterSignal_MASTER/ADDR/$1I2602/I0 ;
  wire \NlwInverterSignal_MASTER/DR_BUS/$1I2913/I0 ;
  wire \NlwInverterSignal_MASTER/DR_BUS/$1I2913/I1 ;
  wire \NlwInverterSignal_MASTER/DR_BUS/$1I2913/I2 ;
  wire \NlwInverterSignal_MASTER/DR_BUS/$1I2805/I0 ;
  wire \NlwInverterSignal_MASTER/DR_BUS/$1I2805/I1 ;
  wire \NlwInverterSignal_MASTER/DR_BUS/$1I2787/I0 ;
  wire \NlwInverterSignal_MASTER/DR_BUS/$1I2752/I0 ;
  wire \NlwInverterSignal_MASTER/DR_BUS/$1I2752/I1 ;
  wire \NlwInverterSignal_MASTER/DR_BUS/$1I2732/I0 ;
  wire \NlwInverterSignal_MASTER/DR_BUS/$1I2732/I1 ;
  wire \NlwInverterSignal_MASTER/DR_BUS/$1I2721/I0 ;
  wire \NlwInverterSignal_MASTER/DR_BUS/$1I2719/I0 ;
  wire \NlwInverterSignal_MASTER/DR_BUS/$1I2706/I0 ;
  wire \NlwInverterSignal_MASTER/DR_BUS/$1I2704/I0 ;
  wire \NlwInverterSignal_MASTER/DR_BUS/$1I2908/$1I7/I0 ;
  wire \NlwInverterSignal_MASTER/DR_BUS/$1I2917/$1I7/I0 ;
  wire \NlwInverterSignal_MASTER/M_DATA/$1I2590/I0 ;
  wire \NlwInverterSignal_MASTER/M_DATA/$1I2518/I0 ;
  wire \NlwInverterSignal_MASTER/M_DATA/$1I2502/I0 ;
  wire \NlwInverterSignal_MASTER/$1I2914/$1I2947/I0 ;
  wire \NlwInverterSignal_MASTER/$1I2914/$1I2931/I0 ;
  wire \NlwInverterSignal_MASTER/$1I2914/$1I2927/I0 ;
  wire \NlwInverterSignal_MASTER/$1I2914/$1I2908/I0 ;
  wire \NlwInverterSignal_MASTER/$1I2914/$1I2895/I0 ;
  wire \NlwInverterSignal_MASTER/$1I2914/$1I2880/I0 ;
  wire \NlwInverterSignal_MASTER/$1I2914/$1I2879/I0 ;
  wire \NlwInverterSignal_MASTER/$1I2914/$1I2853/$1I2213/I0 ;
  wire \NlwInverterSignal_MASTER/$1I2914/$1I2864/$1I2213/I0 ;
  wire \NlwInverterSignal_MASTER/$1I2914/$1I2932/$1I2213/I0 ;
  wire \NlwInverterSignal_MASTER/FRAME/$2I3528/I0 ;
  wire \NlwInverterSignal_MASTER/FRAME/$2I3511/I0 ;
  wire \NlwInverterSignal_MASTER/FRAME/$2I3464/I0 ;
  wire \NlwInverterSignal_MASTER/FRAME/$2I3463/I0 ;
  wire \NlwInverterSignal_MASTER/FRAME/$1I3470/O ;
  wire \NlwInverterSignal_MASTER/FRAME/$1I3466/I0 ;
  wire \NlwInverterSignal_MASTER/FRAME/$1I3393/I0 ;
  wire \NlwInverterSignal_MASTER/FRAME/$1I3368/O ;
  wire \NlwInverterSignal_MASTER/FRAME/$1I3323/I0 ;
  wire \NlwInverterSignal_MASTER/FRAME/$1I3323/O ;
  wire \NlwInverterSignal_MASTER/FRAME/$1I3322/I0 ;
  wire \NlwInverterSignal_MASTER/FRAME/$1I3144/I0 ;
  wire \NlwInverterSignal_MASTER/FRAME/$1I3144/I1 ;
  wire \NlwInverterSignal_MASTER/FRAME/$1I3144/I2 ;
  wire \NLW_MASTER/FRAME/$1I2554/NC_O_UNCONNECTED ;
  wire \NlwInverterSignal_MASTER/FRAME/$1I3467/$1I7/I0 ;
  wire \NlwInverterSignal_MASTER/FRAME/$2I3559/$1I7/I0 ;
  wire \NlwInverterSignal_MASTER/IRDY/$2I3437/I0 ;
  wire \NlwInverterSignal_MASTER/IRDY/$2I3435/O ;
  wire \NlwInverterSignal_MASTER/IRDY/$2I3390/O ;
  wire \NlwInverterSignal_MASTER/IRDY/$2I3332/I0 ;
  wire \NlwInverterSignal_MASTER/IRDY/$2I3332/O ;
  wire \NlwInverterSignal_MASTER/IRDY/$2I3233/I0 ;
  wire \NlwInverterSignal_MASTER/IRDY/$1I3779/I0 ;
  wire \NlwInverterSignal_MASTER/IRDY/$1I3779/O ;
  wire \NlwInverterSignal_MASTER/IRDY/$1I3738/I0 ;
  wire \NlwInverterSignal_MASTER/IRDY/$1I3738/I1 ;
  wire \NlwInverterSignal_MASTER/IRDY/$1I3699/I0 ;
  wire \NlwInverterSignal_MASTER/IRDY/$1I3698/I0 ;
  wire \NlwInverterSignal_MASTER/IRDY/$1I3498/I0 ;
  wire \NlwInverterSignal_MASTER/IRDY/$1I3491/I0 ;
  wire \NlwInverterSignal_MASTER/IRDY/$1I3487/I0 ;
  wire \NlwInverterSignal_MASTER/IRDY/$1I3487/O ;
  wire \NlwInverterSignal_MASTER/IRDY/$1I3211/O ;
  wire \NlwInverterSignal_MASTER/IRDY/$1I3227/$1I7/I0 ;
  wire \NlwInverterSignal_MASTER/IRDY/$1I3492/$1I7/I0 ;
  wire \NlwInverterSignal_MASTER/IRDY/$2I3285/$1I7/I0 ;
  wire \NlwInverterSignal_MASTER/REQ/$1I2726/O ;
  wire \NlwInverterSignal_MASTER/REQ/$1I2721/O ;
  wire \NlwInverterSignal_MASTER/REQ/$1I2670/I0 ;
  wire \NlwInverterSignal_MASTER/REQ/$1I2708/$1I2213/I0 ;
  wire \NlwInverterSignal_MASTER/REQ64/$2I3431/I0 ;
  wire \NlwInverterSignal_MASTER/REQ64/$2I3411/I0 ;
  wire \NlwInverterSignal_MASTER/REQ64/$2I3406/I0 ;
  wire \NlwInverterSignal_MASTER/REQ64/$2I3393/I0 ;
  wire \NlwInverterSignal_MASTER/REQ64/$1I3616/I0 ;
  wire \NlwInverterSignal_MASTER/REQ64/$1I3614/I0 ;
  wire \NlwInverterSignal_MASTER/REQ64/$1I3607/I0 ;
  wire \NlwInverterSignal_MASTER/REQ64/$1I3607/I1 ;
  wire \NlwInverterSignal_MASTER/REQ64/$1I3607/I2 ;
  wire \NlwInverterSignal_MASTER/REQ64/$1I3569/O ;
  wire \NlwInverterSignal_MASTER/REQ64/$1I3561/O ;
  wire \NlwInverterSignal_MASTER/REQ64/$1I3540/I0 ;
  wire \NlwInverterSignal_MASTER/REQ64/$1I3534/I0 ;
  wire \NlwInverterSignal_MASTER/REQ64/$1I3534/O ;
  wire \NLW_MASTER/REQ64/$1I3509/NC_O_UNCONNECTED ;
  wire \NlwInverterSignal_MASTER/REQ64/$1I3562/$1I7/I0 ;
  wire \NlwInverterSignal_MASTER/REQ64/$2I3446/$1I7/I0 ;
  wire \NlwInverterSignal_MASTER/XFERFAIL/$1I3024/I0 ;
  wire \NlwInverterSignal_MASTER/XFERFAIL/$1I3019/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$8I4093/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$8I4047/O ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$8I4045/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$8I4045/I1 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$8I4044/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$8I4044/I1 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$8I4043/O ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$8I4007/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$8I3975/O ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$8I3974/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$8I3974/I1 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$8I3973/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$8I3973/I1 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$8I3971/O ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$7I3977/O ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$7I3976/O ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$7I3975/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$7I3975/I1 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$7I3968/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$7I3968/I1 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$7I3966/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$7I3966/I1 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$7I3965/O ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$6I3740/O ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$6I3739/O ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$6I3738/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$6I3738/I1 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$6I3731/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$6I3731/I1 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$6I3729/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$6I3729/I1 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$6I3728/O ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$5I3899/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$5I3899/O ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$5I3898/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$5I3898/I1 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$5I3898/O ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$5I3893/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$5I3893/O ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$5I3891/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$5I3891/O ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$5I3890/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$5I3890/O ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$5I3889/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$5I3889/O ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$5I3888/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$5I3888/O ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$5I3887/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$5I3887/O ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$5I3886/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$5I3886/O ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$5I3885/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$5I3885/O ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$5I3884/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$5I3884/O ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$5I3883/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$5I3883/I1 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$5I3883/O ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$5I3882/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$5I3882/I1 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$5I3882/O ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$5I3881/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$5I3881/I1 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$5I3881/O ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$4I3785/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$4I3785/O ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$4I3784/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$4I3784/O ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$4I3783/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$4I3783/O ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$4I3782/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$4I3782/O ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$4I3781/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$4I3781/O ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$4I3780/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$4I3780/O ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$4I3779/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$4I3779/I1 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$4I3779/O ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$4I3778/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$4I3778/O ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$4I3776/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$4I3776/O ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$4I3774/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$4I3774/O ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$4I3772/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$4I3772/O ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$4I3770/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$4I3770/I1 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$4I3770/O ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$4I3769/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$4I3769/I1 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$4I3769/O ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$4I3768/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$4I3768/I1 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$4I3768/O ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$3I3105/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$3I3105/I1 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$3I3105/I2 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$3I3105/O ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$3I3093/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$3I3093/I1 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$3I3093/I2 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$3I3093/O ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$2I3723/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$2I3711/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$5I4044/$1I7/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$5I4044/$1I7/I1 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$5I4045/$1I7/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$5I4045/$1I7/I1 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$5I4046/$1I7/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$5I4046/$1I7/I1 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$5I4047/$1I7/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$5I4047/$1I7/I1 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$5I4048/$1I7/I0 ;
  wire \NlwInverterSignal_MASTER/OE_FRAME/$5I4048/$1I7/I1 ;
  wire \NlwInverterSignal_MASTER/S_TAR/$1I2605/I0 ;
  wire \NlwInverterSignal_MASTER/DEV_TO/$1I2789/I0 ;
  wire \NlwInverterSignal_MASTER/DEV_TO/$1I2816/$1I2213/I0 ;
  wire \NlwInverterSignal_MASTER/DEV_TO/$1I2838/$1I2213/I0 ;
  wire \NLW_MASTER/$4I3125/NC_O_UNCONNECTED ;
  wire \NLW_MASTER/$4I3126/NC_O_UNCONNECTED ;
  wire \NLW_MASTER/$4I3127/NC_O_UNCONNECTED ;
  wire \NLW_MASTER/$4I3128/NC_O_UNCONNECTED ;
  wire \NLW_MASTER/$4I3129/NC_O_UNCONNECTED ;
  wire \NLW_MASTER/$4I3130/NC_O_UNCONNECTED ;
  wire \NLW_MASTER/$4I3131/NC_O_UNCONNECTED ;
  wire \NLW_MASTER/$4I3132/NC_O_UNCONNECTED ;
  wire \NLW_MASTER/$4I3134/NC_O_UNCONNECTED ;
  wire \NLW_MASTER/$4I3169/NC_O_UNCONNECTED ;
  wire \NlwInverterSignal_MASTER/LAT_TIMR/$2I56/I0 ;
  wire \NlwInverterSignal_MASTER/LAT_TIMR/$2I56/I1 ;
  wire \NlwInverterSignal_MASTER/LAT_TIMR/$2I56/I2 ;
  wire \NlwInverterSignal_MASTER/LAT_TIMR/$2I23/I0 ;
  wire \NlwInverterSignal_MASTER/LAT_TIMR/$2I23/I1 ;
  wire \NlwInverterSignal_MASTER/LAT_TIMR/$2I23/I2 ;
  wire \NlwInverterSignal_MASTER/LAT_TIMR/$2I23/I3 ;
  wire \NlwInverterSignal_MASTER/LAT_TIMR/$2I21/I0 ;
  wire \NlwInverterSignal_MASTER/LAT_TIMR/$2I21/I1 ;
  wire \NlwInverterSignal_MASTER/LAT_TIMR/$2I21/I2 ;
  wire \NlwInverterSignal_MASTER/LAT_TIMR/$2I19/I0 ;
  wire \NlwInverterSignal_MASTER/LAT_TIMR/$2I19/I1 ;
  wire \NlwInverterSignal_MASTER/LAT_TIMR/$1I8/I0 ;
  wire \NlwInverterSignal_MASTER/LAT_TIMR/$1I8/I1 ;
  wire \NlwInverterSignal_MASTER/LAT_TIMR/$1I29/I0 ;
  wire \NlwInverterSignal_MASTER/LAT_TIMR/$1I29/I1 ;
  wire \NlwInverterSignal_MASTER/LAT_TIMR/$1I29/I2 ;
  wire \NlwInverterSignal_MASTER/LAT_TIMR/$1I29/I3 ;
  wire \NlwInverterSignal_MASTER/LAT_TIMR/$1I25/I0 ;
  wire \NlwInverterSignal_MASTER/LAT_TIMR/$1I25/I1 ;
  wire \NlwInverterSignal_MASTER/LAT_TIMR/$1I25/I2 ;
  wire \NlwInverterSignal_MASTER/LAT_TIMR/$1I11/I0 ;
  wire \NlwInverterSignal_MASTER/LAT_TIMR/Q4/$1I30/$1I7/I0 ;
  wire \NlwInverterSignal_MASTER/LAT_TIMR/Q6/$1I30/$1I7/I0 ;
  wire \NlwInverterSignal_MASTER/LAT_TIMR/Q7/$1I30/$1I7/I0 ;
  wire \NlwInverterSignal_MASTER/LAT_TIMR/TIME_OUT/$1I2214/I0 ;
  wire \NlwInverterSignal_MASTER/LAT_TIMR/Q5/$1I30/$1I7/I0 ;
  wire \NlwInverterSignal_MASTER/LAT_TIMR/Q1/$1I30/$1I7/I0 ;
  wire \NlwInverterSignal_MASTER/LAT_TIMR/Q0/$1I30/$1I7/I0 ;
  wire \NlwInverterSignal_MASTER/LAT_TIMR/Q2/$1I30/$1I7/I0 ;
  wire \NlwInverterSignal_MASTER/LAT_TIMR/Q3/$1I30/$1I7/I0 ;
  wire \NLW_MASTER/PCI-0CH/$1I2529/NC_O_UNCONNECTED ;
  wire \NLW_MASTER/PCI-0CH/$1I2532/NC_O_UNCONNECTED ;
  wire \NLW_MASTER/PCI-0CH/$1I2534/NC_O_UNCONNECTED ;
  wire \NLW_MASTER/PCI-0CH/$1I2536/NC_O_UNCONNECTED ;
  wire \NLW_MASTER/PCI-0CH/$1I2538/NC_O_UNCONNECTED ;
  wire \NLW_MASTER/PCI-0CH/$1I2540/NC_O_UNCONNECTED ;
  wire \NLW_MASTER/PCI-0CH/$1I2542/NC_O_UNCONNECTED ;
  wire \NLW_MASTER/PCI-0CH/$1I2544/NC_O_UNCONNECTED ;
  wire \NLW_MASTER/PCI-0CH/$1I2546/NC_O_UNCONNECTED ;
  wire \NLW_MASTER/PCI-0CH/$1I2548/NC_O_UNCONNECTED ;
  wire \NLW_MASTER/PCI-0CH/$1I2550/NC_O_UNCONNECTED ;
  wire \NLW_MASTER/PCI-0CH/$1I2552/NC_O_UNCONNECTED ;
  wire \NLW_MASTER/PCI-0CH/$1I2554/NC_O_UNCONNECTED ;
  wire \NLW_MASTER/PCI-0CH/$1I2556/NC_O_UNCONNECTED ;
  wire \NLW_MASTER/PCI-0CH/$1I2558/NC_O_UNCONNECTED ;
  wire \NLW_MASTER/PCI-0CH/$1I2560/NC_O_UNCONNECTED ;
  wire \NLW_MASTER/PCI-0CH/$1I2562/NC_O_UNCONNECTED ;
  wire \NLW_MASTER/PCI-0CH/$1I2564/NC_O_UNCONNECTED ;
  wire \NLW_MASTER/PCI-0CH/$1I2566/NC_O_UNCONNECTED ;
  wire \NLW_MASTER/PCI-0CH/$1I2568/NC_O_UNCONNECTED ;
  wire \NLW_MASTER/PCI-0CH/$1I2570/NC_O_UNCONNECTED ;
  wire \NLW_MASTER/PCI-0CH/$1I2572/NC_O_UNCONNECTED ;
  wire \NLW_MASTER/PCI-0CH/$1I2574/NC_O_UNCONNECTED ;
  wire \NLW_MASTER/PCI-0CH/$1I2576/NC_O_UNCONNECTED ;
  wire \NLW_MASTER/PCI-0CH/$1I2578/NC_O_UNCONNECTED ;
  wire \NLW_MASTER/PCI-0CH/$1I2580/NC_O_UNCONNECTED ;
  wire \NLW_MASTER/PCI-0CH/$1I2582/NC_O_UNCONNECTED ;
  wire \NlwInverterSignal_MASTER/3/UPPER/T0/T ;
  wire \NlwInverterSignal_MASTER/3/UPPER/T1/T ;
  wire \NlwInverterSignal_MASTER/3/UPPER/T2/T ;
  wire \NlwInverterSignal_MASTER/3/UPPER/T3/T ;
  wire \NlwInverterSignal_MASTER/3/UPPER/T4/T ;
  wire \NlwInverterSignal_MASTER/3/UPPER/T5/T ;
  wire \NlwInverterSignal_MASTER/3/UPPER/T6/T ;
  wire \NlwInverterSignal_MASTER/3/UPPER/T7/T ;
  wire \NlwInverterSignal_MASTER/3/UPPER/T8/T ;
  wire \NlwInverterSignal_MASTER/3/UPPER/T9/T ;
  wire \NlwInverterSignal_MASTER/3/UPPER/T10/T ;
  wire \NlwInverterSignal_MASTER/3/UPPER/T11/T ;
  wire \NlwInverterSignal_MASTER/3/UPPER/T12/T ;
  wire \NlwInverterSignal_MASTER/3/UPPER/T13/T ;
  wire \NlwInverterSignal_MASTER/3/UPPER/T14/T ;
  wire \NlwInverterSignal_MASTER/3/UPPER/T15/T ;
  wire \NlwInverterSignal_MASTER/3/LOWER/T0/T ;
  wire \NlwInverterSignal_MASTER/3/LOWER/T1/T ;
  wire \NlwInverterSignal_MASTER/3/LOWER/T2/T ;
  wire \NlwInverterSignal_MASTER/3/LOWER/T3/T ;
  wire \NlwInverterSignal_MASTER/3/LOWER/T4/T ;
  wire \NlwInverterSignal_MASTER/3/LOWER/T5/T ;
  wire \NlwInverterSignal_MASTER/3/LOWER/T6/T ;
  wire \NlwInverterSignal_MASTER/3/LOWER/T7/T ;
  wire \NlwInverterSignal_MASTER/3/LOWER/T8/T ;
  wire \NlwInverterSignal_MASTER/3/LOWER/T9/T ;
  wire \NlwInverterSignal_MASTER/3/LOWER/T10/T ;
  wire \NlwInverterSignal_MASTER/3/LOWER/T11/T ;
  wire \NlwInverterSignal_MASTER/3/LOWER/T12/T ;
  wire \NlwInverterSignal_MASTER/3/LOWER/T13/T ;
  wire \NlwInverterSignal_MASTER/3/LOWER/T14/T ;
  wire \NlwInverterSignal_MASTER/3/LOWER/T15/T ;
  wire \NLW_MASTER/$4I3247/NC_O_UNCONNECTED ;
  wire \NLW_MASTER/$4I3298/NC_O_UNCONNECTED ;
  wire \NLW_MASTER/$4I3318/NC_O_UNCONNECTED ;
  wire \NlwInverterSignal_PCI-CNTL/$4I788/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/$4I719/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/$4I446/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/$1I840/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/$1I840/I1 ;
  wire \NlwInverterSignal_PCI-CNTL/$1I823/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/$1I1005/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-LC/$2I3201/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-LC/$2I3201/I1 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-LC/$2I3192/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-LC/$2I3076/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OE/$2I940/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OE/$2I934/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OE/$2I933/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OE/$2I932/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OE/$2I777/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OE/$2I777/I1 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OE/$2I592/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OE/OE15/$1I307/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OE/OE15/$1I296/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OE/OE7/$1I307/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OE/OE7/$1I296/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OE/OE6/$1I307/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OE/OE6/$1I296/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OE/OE5/$1I307/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OE/OE5/$1I296/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OE/OE4/$1I307/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OE/OE4/$1I296/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OE/OE3/$1I307/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OE/OE3/$1I296/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OE/OE8/$1I307/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OE/OE8/$1I296/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OE/OE9/$1I307/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OE/OE9/$1I296/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OE/OE12/$1I307/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OE/OE12/$1I296/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OE/OE1/$1I307/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OE/OE1/$1I296/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OE/$2I617/$1I11/I0 ;
  wire \NLW_PCI-CNTL/PCI-OE/SW1/$1I2289/NC_O_UNCONNECTED ;
  wire \NLW_PCI-CNTL/PCI-OE/SW15/$1I2289/NC_O_UNCONNECTED ;
  wire \NLW_PCI-CNTL/PCI-OE/SW3/$1I2289/NC_O_UNCONNECTED ;
  wire \NLW_PCI-CNTL/$1I972/NC_O_UNCONNECTED ;
  wire \NLW_PCI-CNTL/$1I974/NC_O_UNCONNECTED ;
  wire \NlwInverterSignal_PCI-CNTL/$1I995/$1I2213/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-IDLE/$1I494/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-IDLE/$1I494/I1 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-BUSY/$1I542/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-BUSY/$1I521/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-BUSY/$1I471/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-BUSY/$1I471/I1 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-BUSY/$1I469/I0 ;
  wire \NLW_PCI-CNTL/PCI-TSM/PCI-BUSY/$1I587/NC_O_UNCONNECTED ;
  wire \NLW_PCI-CNTL/PCI-TSM/PCI-BUSY/$1I588/NC_O_UNCONNECTED ;
  wire \NLW_PCI-CNTL/PCI-TSM/PCI-BUSY/$1I589/NC_O_UNCONNECTED ;
  wire \NLW_PCI-CNTL/PCI-TSM/PCI-BUSY/$1I590/NC_O_UNCONNECTED ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-DATA/$1I670/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-DATA/$1I670/I1 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-DATA/$1I627/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-DATA/$1I481/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-DATA/$1I480/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-DATA/$1I480/I1 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-DATA/$1I480/I2 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-DATA/$1I453/I0 ;
  wire \NLW_PCI-CNTL/PCI-TSM/PCI-DATA/$1I568/NC_O_UNCONNECTED ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-BKOF/$1I579/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-BKOF/$1I575/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-BKOF/$1I526/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-BKOF/$1I526/I1 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-BKOF/$1I486/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-BKOF/$1I475/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-BKOF/$1I474/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-BKOF/$1I474/I1 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-BKOF/$1I458/I0 ;
  wire \NLW_PCI-CNTL/PCI-TSM/$1I489/NC_O_UNCONNECTED ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-AK64/$3I855/O ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-AK64/$2I971/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-AK64/$2I965/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-AK64/$2I958/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-AK64/$2I951/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-AK64/$2I941/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-AK64/$1I837/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-AK64/$1I797/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-AK64/$1I796/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-AK64/$1I787/O ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-AK64/$1I781/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-AK64/$1I781/I1 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-AK64/$3I854/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-DSEL/$3I795/O ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-DSEL/$2I983/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-DSEL/$2I951/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-DSEL/$2I931/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-DSEL/$2I914/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-DSEL/$2I878/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-DSEL/$1I801/O ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-DSEL/$1I768/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-DSEL/$1I760/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-DSEL/$1I758/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-DSEL/$1I1028/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-DSEL/$1I1028/I1 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-DSEL/$3I798/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$4I977/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$4I1044/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$4I1044/I1 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$4I1010/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$4I1010/O ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$3I856/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$3I856/I1 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$3I825/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$3I823/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$3I822/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$3I616/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$3I616/O ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I785/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I768/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I746/O ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I731/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I481/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I480/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I480/I1 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I480/I2 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I459/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I459/I1 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I453/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I782/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$4I1028/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$3I1287/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$3I1287/O ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$3I1286/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$3I1284/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$3I1263/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$3I1263/O ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$3I1260/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$3I1258/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1504/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1480/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1450/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1248/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1060/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1368/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1373/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1437/$1I2213/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1499/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$6I970/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$6I970/O ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$6I969/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$6I969/O ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$6I966/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$6I966/O ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$6I965/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$6I965/O ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$5I1041/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$5I1035/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$5I1035/I1 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$5I1034/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$5I1034/I1 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$4I909/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$4I909/O ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$4I908/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$4I908/O ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$4I905/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$4I905/O ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$4I903/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$4I903/O ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$3I899/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$3I890/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$3I890/I1 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$3I801/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$3I801/I1 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$3I627/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$2I822/O ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$2I1330/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$2I1330/I1 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$2I1330/I2 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$2I1265/O ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$2I1014/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$2I1014/I1 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$2I1014/I2 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$1I1251/I0 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$1I1251/I1 ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$1I1251/O ;
  wire \NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$1I1247/I0 ;
  wire \NLW_PCI-CNTL/PCI-OFCN/PCI-XOE/$1I1031/NC_O_UNCONNECTED ;
  wire \NLW_PCI-CNTL/PCI-OFCN/PCI-XOE/$1I1065/NC_O_UNCONNECTED ;
  wire \NLW_PCI-CNTL/PCI-OFCN/PCI-XOE/$1I1239/NC_O_UNCONNECTED ;
  wire \NLW_PCI-CNTL/PCI-OFCN/PCI-XOE/$1I1240/NC_O_UNCONNECTED ;
  wire \NLW_PCI-CNTL/$3I992/NC_O_UNCONNECTED ;
  wire \NlwInverterSignal_PCI-CNTL/$4I614/$1I7/I0 ;
  wire \NLW_$1I3754/NC_O_UNCONNECTED ;
  wire \NLW_$1I3755/NC_O_UNCONNECTED ;
  wire \NLW_$1I3756/NC_O_UNCONNECTED ;
  wire \NLW_$1I3757/NC_O_UNCONNECTED ;
  wire \NLW_$1I3758/NC_O_UNCONNECTED ;
  wire \NLW_$1I3759/NC_O_UNCONNECTED ;
  wire \NLW_$1I3760/NC_O_UNCONNECTED ;
  wire \NLW_$1I3761/NC_O_UNCONNECTED ;
  wire \NLW_$1I3762/NC_O_UNCONNECTED ;
  wire \NLW_$1I3763/NC_O_UNCONNECTED ;
  wire \NLW_$1I3764/NC_O_UNCONNECTED ;
  wire \NLW_$1I3765/NC_O_UNCONNECTED ;
  wire \NLW_$1I3766/NC_O_UNCONNECTED ;
  wire \NLW_$1I3767/NC_O_UNCONNECTED ;
  wire \NLW_$1I3768/NC_O_UNCONNECTED ;
  wire \NLW_$1I3769/NC_O_UNCONNECTED ;
  wire \NLW_$1I3770/NC_O_UNCONNECTED ;
  wire \NLW_$1I3771/NC_O_UNCONNECTED ;
  wire \NLW_$1I3772/NC_O_UNCONNECTED ;
  wire \NLW_$1I3773/NC_O_UNCONNECTED ;
  wire \NLW_$1I3774/NC_O_UNCONNECTED ;
  wire \NLW_$1I3775/NC_O_UNCONNECTED ;
  wire \NLW_$1I3776/NC_O_UNCONNECTED ;
  wire \NLW_$1I3777/NC_O_UNCONNECTED ;
  wire \NLW_$1I3778/NC_O_UNCONNECTED ;
  wire \NLW_$1I3779/NC_O_UNCONNECTED ;
  wire \NLW_$1I3780/NC_O_UNCONNECTED ;
  wire \NLW_$1I3781/NC_O_UNCONNECTED ;
  wire \NLW_$1I3782/NC_O_UNCONNECTED ;
  wire \NLW_$1I3783/NC_O_UNCONNECTED ;
  wire \NLW_$1I3784/NC_O_UNCONNECTED ;
  wire \NLW_$1I3785/NC_O_UNCONNECTED ;
  wire \NLW_$1I3786/NC_O_UNCONNECTED ;
  wire \NLW_$1I3787/NC_O_UNCONNECTED ;
  wire \NLW_$1I3788/NC_O_UNCONNECTED ;
  wire \NLW_$1I3789/NC_O_UNCONNECTED ;
  wire \NLW_$1I3790/NC_O_UNCONNECTED ;
  wire \NLW_$1I3791/NC_O_UNCONNECTED ;
  wire \NLW_$1I3792/NC_O_UNCONNECTED ;
  wire \NLW_$1I3793/NC_O_UNCONNECTED ;
  wire \NLW_$1I3794/NC_O_UNCONNECTED ;
  wire \NLW_$1I3795/NC_O_UNCONNECTED ;
  wire \NLW_$1I3796/NC_O_UNCONNECTED ;
  wire \NLW_$1I3797/NC_O_UNCONNECTED ;
  wire \NLW_$1I3798/NC_O_UNCONNECTED ;
  wire \NLW_$1I3799/NC_O_UNCONNECTED ;
  wire \NLW_$1I3800/NC_O_UNCONNECTED ;
  wire \NLW_$1I3801/NC_O_UNCONNECTED ;
  wire \NLW_$1I3802/NC_O_UNCONNECTED ;
  wire \NLW_$1I3803/NC_O_UNCONNECTED ;
  wire \NLW_$1I3804/NC_O_UNCONNECTED ;
  wire \NLW_$1I3805/NC_O_UNCONNECTED ;
  wire \NLW_$1I3806/NC_O_UNCONNECTED ;
  wire \NLW_$1I3807/NC_O_UNCONNECTED ;
  wire \NLW_$1I3808/NC_O_UNCONNECTED ;
  wire \NLW_$1I3809/NC_O_UNCONNECTED ;
  wire \NLW_$1I3810/NC_O_UNCONNECTED ;
  wire \NLW_$1I3811/NC_O_UNCONNECTED ;
  wire \NLW_$1I3812/NC_O_UNCONNECTED ;
  wire \NLW_$1I3813/NC_O_UNCONNECTED ;
  wire \NLW_$1I3814/NC_O_UNCONNECTED ;
  wire \NLW_$1I3815/NC_O_UNCONNECTED ;
  wire \NLW_$1I3816/NC_O_UNCONNECTED ;
  wire \NLW_$1I3817/NC_O_UNCONNECTED ;
  wire \NLW_$1I3818/NC_O_UNCONNECTED ;
  wire \NLW_$1I3819/NC_O_UNCONNECTED ;
  wire \NLW_$1I3820/NC_O_UNCONNECTED ;
  wire \NLW_$1I3821/NC_O_UNCONNECTED ;
  wire \NLW_$1I3822/NC_O_UNCONNECTED ;
  wire \NLW_$1I3823/NC_O_UNCONNECTED ;
  wire \NLW_$1I3824/NC_O_UNCONNECTED ;
  wire \NLW_$1I3825/NC_O_UNCONNECTED ;
  wire \NLW_$1I3826/NC_O_UNCONNECTED ;
  wire \NLW_$1I3827/NC_O_UNCONNECTED ;
  wire \NLW_$1I3828/NC_O_UNCONNECTED ;
  wire \NLW_$1I3829/NC_O_UNCONNECTED ;
  wire \NLW_$1I3830/NC_O_UNCONNECTED ;
  wire \NLW_$1I3831/NC_O_UNCONNECTED ;
  wire \NLW_$1I3832/NC_O_UNCONNECTED ;
  wire \NLW_$1I3833/NC_O_UNCONNECTED ;
  wire \NLW_$1I3834/NC_O_UNCONNECTED ;
  wire \NLW_$1I3835/NC_O_UNCONNECTED ;
  wire \NLW_$1I3836/NC_O_UNCONNECTED ;
  wire \NLW_$1I3837/NC_O_UNCONNECTED ;
  wire \NLW_$1I3840/NC_O_UNCONNECTED ;
  wire \NLW_$1I3841/NC_O_UNCONNECTED ;
  wire \NLW_$1I3842/NC_O_UNCONNECTED ;
  wire \NLW_$1I3843/NC_O_UNCONNECTED ;
  wire \NLW_$1I3844/NC_O_UNCONNECTED ;
  wire \NLW_$1I3845/NC_O_UNCONNECTED ;
  wire \NLW_$1I3846/NC_O_UNCONNECTED ;
  wire \NLW_$1I3847/NC_O_UNCONNECTED ;
  wire \NLW_$1I3848/NC_O_UNCONNECTED ;
  wire \NLW_$1I3849/NC_O_UNCONNECTED ;
  wire \NLW_$1I3850/NC_O_UNCONNECTED ;
  wire \NLW_$1I3851/NC_O_UNCONNECTED ;
  wire \NLW_$1I3852/NC_O_UNCONNECTED ;
  wire \NLW_$1I3853/NC_O_UNCONNECTED ;
  wire \NLW_$1I3854/NC_O_UNCONNECTED ;
  wire \NLW_$1I3855/NC_O_UNCONNECTED ;
  wire \NLW_$1I3860/NC_O_UNCONNECTED ;
  wire \NLW_$1I3861/NC_O_UNCONNECTED ;
  wire \NLW_$1I3862/NC_O_UNCONNECTED ;
  wire \NLW_$1I3863/NC_O_UNCONNECTED ;
  wire \NLW_$1I3864/NC_O_UNCONNECTED ;
  wire \NLW_$1I3865/NC_O_UNCONNECTED ;
  wire \NLW_$1I3866/NC_O_UNCONNECTED ;
  wire \NLW_$1I3867/NC_O_UNCONNECTED ;
  wire \NLW_$1I3868/NC_O_UNCONNECTED ;
  wire \NLW_$1I3869/NC_O_UNCONNECTED ;
  wire \NLW_$1I3870/NC_O_UNCONNECTED ;
  wire \NLW_$1I3871/NC_O_UNCONNECTED ;
  wire \NLW_$1I3872/NC_O_UNCONNECTED ;
  wire \NLW_$1I3873/NC_O_UNCONNECTED ;
  wire \NLW_$1I3874/NC_O_UNCONNECTED ;
  wire \NLW_$1I3875/NC_O_UNCONNECTED ;
  wire \NLW_$1I3879/NC_O_UNCONNECTED ;
  wire \NLW_$1I3880/NC_O_UNCONNECTED ;
  wire \NLW_$1I3881/NC_O_UNCONNECTED ;
  wire \NLW_$1I3882/NC_O_UNCONNECTED ;
  wire \NLW_$1I3883/NC_O_UNCONNECTED ;
  wire \NLW_$1I3884/NC_O_UNCONNECTED ;
  wire \NLW_$1I3885/NC_O_UNCONNECTED ;
  wire \NLW_$1I3886/NC_O_UNCONNECTED ;
  wire \NLW_$1I3887/NC_O_UNCONNECTED ;
  wire \NLW_$1I3888/NC_O_UNCONNECTED ;
  wire \NLW_$1I3889/NC_O_UNCONNECTED ;
  wire \NLW_$1I3890/NC_O_UNCONNECTED ;
  wire \NLW_$1I3891/NC_O_UNCONNECTED ;
  wire \NLW_$1I3892/NC_O_UNCONNECTED ;
  wire \NLW_$1I3893/NC_O_UNCONNECTED ;
  wire \NLW_$1I3894/NC_O_UNCONNECTED ;
  wire \NLW_$1I3895/NC_O_UNCONNECTED ;
  wire \NLW_$1I3896/NC_O_UNCONNECTED ;
  wire \NLW_$1I3897/NC_O_UNCONNECTED ;
  wire \NLW_$1I3898/NC_O_UNCONNECTED ;
  wire \NLW_$1I3899/NC_O_UNCONNECTED ;
  wire \NLW_$1I3900/NC_O_UNCONNECTED ;
  wire \NLW_$1I3901/NC_O_UNCONNECTED ;
  wire \NLW_$1I3902/NC_O_UNCONNECTED ;
  wire \NLW_$1I3903/NC_O_UNCONNECTED ;
  wire \NLW_$1I3904/NC_O_UNCONNECTED ;
  wire \NLW_$1I3905/NC_O_UNCONNECTED ;
  wire \NLW_$1I3906/NC_O_UNCONNECTED ;
  wire \NLW_$1I3907/NC_O_UNCONNECTED ;
  wire \NLW_$1I3908/NC_O_UNCONNECTED ;
  wire \NLW_$1I3909/NC_O_UNCONNECTED ;
  wire \NLW_$1I3910/NC_O_UNCONNECTED ;
  wire \NLW_$1I3911/NC_O_UNCONNECTED ;
  wire \NLW_$1I3912/NC_O_UNCONNECTED ;
  wire \NLW_$1I3913/NC_O_UNCONNECTED ;
  wire \NLW_$1I3914/NC_O_UNCONNECTED ;
  wire \NLW_$1I3915/NC_O_UNCONNECTED ;
  wire \NLW_$1I3916/NC_O_UNCONNECTED ;
  wire \NLW_$1I3917/NC_O_UNCONNECTED ;
  wire \NLW_$1I3918/NC_O_UNCONNECTED ;
  wire \NLW_$1I3921/NC_O_UNCONNECTED ;
  wire \NLW_$1I3922/NC_O_UNCONNECTED ;
  wire \NLW_$1I3923/NC_O_UNCONNECTED ;
  wire \NLW_$1I3924/NC_O_UNCONNECTED ;
  wire \NLW_$1I3925/NC_O_UNCONNECTED ;
  wire \NLW_$1I3926/NC_O_UNCONNECTED ;
  wire \NLW_$1I3927/NC_O_UNCONNECTED ;
  wire \NLW_$1I3928/NC_O_UNCONNECTED ;
  wire \NLW_$1I4355/NC_O_UNCONNECTED ;
  wire \NLW_$1I4356/NC_O_UNCONNECTED ;
  wire \NLW_$1I4357/NC_O_UNCONNECTED ;
  wire \NLW_$1I4358/NC_O_UNCONNECTED ;
  wire \NLW_$1I4359/NC_O_UNCONNECTED ;
  wire \NLW_$1I4360/NC_O_UNCONNECTED ;
  wire \NLW_$1I4361/NC_O_UNCONNECTED ;
  wire \NLW_$1I4362/NC_O_UNCONNECTED ;
  wire \NLW_$1I4363/NC_O_UNCONNECTED ;
  wire \NLW_$1I4364/NC_O_UNCONNECTED ;
  wire \NLW_$1I4365/NC_O_UNCONNECTED ;
  wire \NLW_$1I4366/NC_O_UNCONNECTED ;
  wire \NLW_$1I4367/NC_O_UNCONNECTED ;
  wire \NLW_$1I4368/NC_O_UNCONNECTED ;
  wire \NLW_$1I4369/NC_O_UNCONNECTED ;
  wire \NLW_$1I4370/NC_O_UNCONNECTED ;
  wire \NLW_$1I4371/NC_O_UNCONNECTED ;
  wire \NLW_$1I4372/NC_O_UNCONNECTED ;
  wire \NLW_$1I4373/NC_O_UNCONNECTED ;
  wire \NLW_$1I4374/NC_O_UNCONNECTED ;
  wire \NLW_$1I4375/NC_O_UNCONNECTED ;
  wire \NLW_$1I4376/NC_O_UNCONNECTED ;
  wire \NLW_$1I4377/NC_O_UNCONNECTED ;
  wire \NLW_$1I4378/NC_O_UNCONNECTED ;
  wire \NLW_$1I4379/NC_O_UNCONNECTED ;
  wire \NLW_$1I4380/NC_O_UNCONNECTED ;
  wire \NLW_$1I4381/NC_O_UNCONNECTED ;
  wire \NLW_$1I4382/NC_O_UNCONNECTED ;
  wire \NLW_$1I4383/NC_O_UNCONNECTED ;
  wire \NLW_$1I4384/NC_O_UNCONNECTED ;
  wire \NLW_$1I4385/NC_O_UNCONNECTED ;
  wire \NLW_$1I4386/NC_O_UNCONNECTED ;
  wire \NLW_$1I4387/NC_O_UNCONNECTED ;
  wire \NLW_$1I4388/NC_O_UNCONNECTED ;
  wire \NLW_$1I4389/NC_O_UNCONNECTED ;
  wire \NLW_$1I4390/NC_O_UNCONNECTED ;
  wire \NLW_$1I4391/NC_O_UNCONNECTED ;
  wire \NLW_$1I4392/NC_O_UNCONNECTED ;
  wire \NLW_$1I4393/NC_O_UNCONNECTED ;
  wire \NLW_$1I4394/NC_O_UNCONNECTED ;
  wire \NLW_$1I4395/NC_O_UNCONNECTED ;
  wire \NLW_$1I4396/NC_O_UNCONNECTED ;
  wire \NLW_$1I4397/NC_O_UNCONNECTED ;
  wire \NLW_$1I4398/NC_O_UNCONNECTED ;
  wire \NLW_$1I4399/NC_O_UNCONNECTED ;
  wire \NLW_$1I4400/NC_O_UNCONNECTED ;
  wire \NLW_$1I4401/NC_O_UNCONNECTED ;
  wire \NLW_$1I4402/NC_O_UNCONNECTED ;
  wire \NLW_$1I4403/NC_O_UNCONNECTED ;
  wire \NLW_$1I4404/NC_O_UNCONNECTED ;
  wire \NLW_$1I4405/NC_O_UNCONNECTED ;
  wire \NLW_$1I4406/NC_O_UNCONNECTED ;
  wire \NLW_$1I4407/NC_O_UNCONNECTED ;
  wire \NLW_$1I4408/NC_O_UNCONNECTED ;
  wire \NLW_$1I4409/NC_O_UNCONNECTED ;
  wire \NLW_$1I4410/NC_O_UNCONNECTED ;
  wire \NLW_$1I4411/NC_O_UNCONNECTED ;
  wire \NLW_$1I4412/NC_O_UNCONNECTED ;
  wire \NLW_$1I4413/NC_O_UNCONNECTED ;
  wire \NLW_$1I4414/NC_O_UNCONNECTED ;
  wire \NLW_$1I4415/NC_O_UNCONNECTED ;
  wire \NLW_$1I4416/NC_O_UNCONNECTED ;
  wire \NLW_$1I4417/NC_O_UNCONNECTED ;
  wire \NLW_$1I4418/NC_O_UNCONNECTED ;
  wire \NLW_$1I4419/NC_O_UNCONNECTED ;
  wire \NLW_$1I4420/NC_O_UNCONNECTED ;
  wire \NLW_$1I4421/NC_O_UNCONNECTED ;
  wire \NLW_$1I4422/NC_O_UNCONNECTED ;
  wire \NLW_$1I4423/NC_O_UNCONNECTED ;
  wire \NLW_$1I4424/NC_O_UNCONNECTED ;
  wire \NLW_$1I4425/NC_O_UNCONNECTED ;
  wire \NLW_$1I4426/NC_O_UNCONNECTED ;
  wire \NLW_$1I4427/NC_O_UNCONNECTED ;
  wire \NLW_$1I4428/NC_O_UNCONNECTED ;
  wire \NLW_$1I4429/NC_O_UNCONNECTED ;
  wire \NLW_$1I4430/NC_O_UNCONNECTED ;
  wire \NLW_$1I4431/NC_O_UNCONNECTED ;
  wire \NLW_$1I4432/NC_O_UNCONNECTED ;
  wire \NLW_$1I4433/NC_O_UNCONNECTED ;
  wire \NLW_$1I4434/NC_O_UNCONNECTED ;
  wire \NLW_$1I4435/NC_O_UNCONNECTED ;
  wire \NLW_$1I4436/NC_O_UNCONNECTED ;
  wire \NLW_$1I4437/NC_O_UNCONNECTED ;
  wire \NLW_$1I4438/NC_O_UNCONNECTED ;
  wire \NLW_$1I4439/NC_O_UNCONNECTED ;
  wire \NLW_$1I4440/NC_O_UNCONNECTED ;
  wire \NLW_$1I4441/NC_O_UNCONNECTED ;
  wire \NLW_$1I4442/NC_O_UNCONNECTED ;
  wire \NLW_$1I4443/NC_O_UNCONNECTED ;
  wire \NLW_$1I4444/NC_O_UNCONNECTED ;
  wire \NLW_$1I4445/NC_O_UNCONNECTED ;
  wire \NLW_$1I4446/NC_O_UNCONNECTED ;
  wire \NLW_$1I4447/NC_O_UNCONNECTED ;
  wire \NLW_$1I4448/NC_O_UNCONNECTED ;
  wire \NLW_$1I4449/NC_O_UNCONNECTED ;
  wire \NLW_$1I4450/NC_O_UNCONNECTED ;
  wire \NLW_$1I4451/NC_O_UNCONNECTED ;
  wire \NLW_$1I4452/NC_O_UNCONNECTED ;
  wire \NLW_$1I4453/NC_O_UNCONNECTED ;
  wire \NLW_$1I4454/NC_O_UNCONNECTED ;
  wire \NLW_$1I4455/NC_O_UNCONNECTED ;
  wire \NLW_$1I4456/NC_O_UNCONNECTED ;
  wire \NLW_$1I4457/NC_O_UNCONNECTED ;
  wire \NLW_$1I4458/NC_O_UNCONNECTED ;
  wire \NLW_$1I4459/NC_O_UNCONNECTED ;
  wire \NLW_$1I4460/NC_O_UNCONNECTED ;
  wire \NLW_$1I4461/NC_O_UNCONNECTED ;
  wire \NLW_$1I4462/NC_O_UNCONNECTED ;
  wire \NLW_$1I4463/NC_O_UNCONNECTED ;
  wire \NLW_$1I4464/NC_O_UNCONNECTED ;
  wire \NLW_$1I4465/NC_O_UNCONNECTED ;
  wire \NLW_$1I4466/NC_O_UNCONNECTED ;
  wire \NLW_$1I4467/NC_O_UNCONNECTED ;
  wire \NLW_$1I4468/NC_O_UNCONNECTED ;
  wire \NLW_$1I4469/NC_O_UNCONNECTED ;
  wire \NLW_$1I4470/NC_O_UNCONNECTED ;
  wire \NLW_$1I4471/NC_O_UNCONNECTED ;
  wire \NLW_$1I4472/NC_O_UNCONNECTED ;
  wire \NLW_$1I4473/NC_O_UNCONNECTED ;
  wire \NLW_$1I4474/NC_O_UNCONNECTED ;
  wire \NLW_$1I4475/NC_O_UNCONNECTED ;
  wire \NLW_$1I4476/NC_O_UNCONNECTED ;
  wire \NLW_$1I4477/NC_O_UNCONNECTED ;
  wire \NLW_$1I4478/NC_O_UNCONNECTED ;
  wire \NLW_$1I4479/NC_O_UNCONNECTED ;
  wire \NLW_$1I4480/NC_O_UNCONNECTED ;
  wire \NLW_$1I4481/NC_O_UNCONNECTED ;
  wire \NLW_$1I4482/NC_O_UNCONNECTED ;
  wire \NLW_$1I4483/NC_O_UNCONNECTED ;
  wire \NLW_$1I4484/NC_O_UNCONNECTED ;
  wire \NLW_$1I4485/NC_O_UNCONNECTED ;
  wire \NLW_$1I4486/NC_O_UNCONNECTED ;
  wire \NLW_$1I4487/NC_O_UNCONNECTED ;
  wire \NLW_$1I4488/NC_O_UNCONNECTED ;
  wire \NLW_$1I4489/NC_O_UNCONNECTED ;
  wire \NLW_$1I4490/NC_O_UNCONNECTED ;
  wire \NLW_$1I4491/NC_O_UNCONNECTED ;
  wire \NLW_$1I4492/NC_O_UNCONNECTED ;
  wire \NLW_$1I4493/NC_O_UNCONNECTED ;
  wire \NLW_$1I4494/NC_O_UNCONNECTED ;
  wire \NLW_$1I4495/NC_O_UNCONNECTED ;
  wire \NLW_$1I4496/NC_O_UNCONNECTED ;
  wire \NLW_$1I4497/NC_O_UNCONNECTED ;
  wire \NLW_$1I4498/NC_O_UNCONNECTED ;
  wire \NLW_$1I4499/NC_O_UNCONNECTED ;
  wire \NLW_$1I4500/NC_O_UNCONNECTED ;
  wire \NLW_$1I4501/NC_O_UNCONNECTED ;
  wire \NLW_$1I4502/NC_O_UNCONNECTED ;
  wire \NLW_$1I4503/NC_O_UNCONNECTED ;
  wire \NLW_$1I4504/NC_O_UNCONNECTED ;
  wire \NLW_$1I4505/NC_O_UNCONNECTED ;
  wire \NLW_$1I4506/NC_O_UNCONNECTED ;
  wire \NLW_$1I4507/NC_O_UNCONNECTED ;
  wire \NLW_$1I4508/NC_O_UNCONNECTED ;
  wire \NLW_$1I4509/NC_O_UNCONNECTED ;
  wire \NLW_$1I4510/NC_O_UNCONNECTED ;
  wire \NLW_$1I4511/NC_O_UNCONNECTED ;
  wire \NLW_$1I4512/NC_O_UNCONNECTED ;
  wire \NLW_$1I4513/NC_O_UNCONNECTED ;
  wire \NLW_$1I4514/NC_O_UNCONNECTED ;
  wire \NLW_$1I4515/NC_O_UNCONNECTED ;
  wire \NLW_$1I4516/NC_O_UNCONNECTED ;
  wire \NLW_$1I4517/NC_O_UNCONNECTED ;
  wire \NLW_$1I4518/NC_O_UNCONNECTED ;
  wire \NLW_$1I4519/NC_O_UNCONNECTED ;
  wire \NLW_$1I4520/NC_O_UNCONNECTED ;
  wire \NLW_$1I4521/NC_O_UNCONNECTED ;
  wire \NLW_$1I4522/NC_O_UNCONNECTED ;
  wire \NLW_$1I4523/NC_O_UNCONNECTED ;
  wire \NLW_$1I4524/NC_O_UNCONNECTED ;
  wire \NLW_$1I4525/NC_O_UNCONNECTED ;
  wire \NLW_$1I4526/NC_O_UNCONNECTED ;
  wire \NLW_$1I4527/NC_O_UNCONNECTED ;
  wire \NLW_$1I4528/NC_O_UNCONNECTED ;
  wire \NLW_$1I4529/NC_O_UNCONNECTED ;
  wire \NLW_$1I4530/NC_O_UNCONNECTED ;
  wire \NLW_$1I4531/NC_O_UNCONNECTED ;
  wire \NLW_$1I4532/NC_O_UNCONNECTED ;
  wire \NLW_$1I4533/NC_O_UNCONNECTED ;
  wire \NLW_$1I4534/NC_O_UNCONNECTED ;
  wire \NLW_$1I4535/NC_O_UNCONNECTED ;
  wire \NLW_$1I4536/NC_O_UNCONNECTED ;
  wire \NLW_$1I4537/NC_O_UNCONNECTED ;
  wire \NLW_$1I4538/NC_O_UNCONNECTED ;
  wire \NLW_$1I4539/NC_O_UNCONNECTED ;
  wire \NLW_$1I4540/NC_O_UNCONNECTED ;
  wire \NLW_$1I4541/NC_O_UNCONNECTED ;
  wire \NLW_$1I4542/NC_O_UNCONNECTED ;
  wire \NLW_$1I4543/NC_O_UNCONNECTED ;
  wire \NLW_$1I4544/NC_O_UNCONNECTED ;
  wire \NLW_$1I4545/NC_O_UNCONNECTED ;
  wire \NLW_$1I4546/NC_O_UNCONNECTED ;
  wire \NLW_$1I4547/NC_O_UNCONNECTED ;
  wire \NLW_$1I4548/NC_O_UNCONNECTED ;
  wire \NLW_$1I4549/NC_O_UNCONNECTED ;
  wire \NLW_$1I4550/NC_O_UNCONNECTED ;
  wire \NLW_$1I4551/NC_O_UNCONNECTED ;
  wire \NLW_$1I4552/NC_O_UNCONNECTED ;
  wire \NLW_$1I4553/NC_O_UNCONNECTED ;
  wire \NLW_$1I4554/NC_O_UNCONNECTED ;
  wire \NLW_$1I4555/NC_O_UNCONNECTED ;
  wire \NLW_$1I4556/NC_O_UNCONNECTED ;
  wire \NLW_$1I4557/NC_O_UNCONNECTED ;
  wire \NLW_$1I4558/NC_O_UNCONNECTED ;
  wire \NLW_$1I4559/NC_O_UNCONNECTED ;
  wire \NLW_$1I4560/NC_O_UNCONNECTED ;
  wire \NLW_$1I4561/NC_O_UNCONNECTED ;
  wire \NLW_$1I4562/NC_O_UNCONNECTED ;
  wire \NLW_$1I4563/NC_O_UNCONNECTED ;
  wire \NLW_$1I4564/NC_O_UNCONNECTED ;
  wire \NLW_$1I4565/NC_O_UNCONNECTED ;
  wire \NLW_$1I4566/NC_O_UNCONNECTED ;
  wire \NLW_$1I4567/NC_O_UNCONNECTED ;
  wire \NLW_$1I4568/NC_O_UNCONNECTED ;
  wire \NLW_$1I4569/NC_O_UNCONNECTED ;
  wire \NLW_$1I4570/NC_O_UNCONNECTED ;
  wire \NLW_$1I4571/NC_O_UNCONNECTED ;
  wire \NLW_$1I4572/NC_O_UNCONNECTED ;
  wire \NLW_$1I4573/NC_O_UNCONNECTED ;
  wire \NLW_$1I4574/NC_O_UNCONNECTED ;
  wire \NLW_$1I4575/NC_O_UNCONNECTED ;
  wire \NLW_$1I4576/NC_O_UNCONNECTED ;
  wire \NLW_$1I4577/NC_O_UNCONNECTED ;
  wire \NLW_$1I4578/NC_O_UNCONNECTED ;
  wire \NLW_$1I4579/NC_O_UNCONNECTED ;
  wire \NLW_$1I4580/NC_O_UNCONNECTED ;
  wire \NLW_$1I4581/NC_O_UNCONNECTED ;
  wire \NLW_$1I4582/NC_O_UNCONNECTED ;
  wire \NLW_$1I4583/NC_O_UNCONNECTED ;
  wire \NLW_$1I4584/NC_O_UNCONNECTED ;
  wire \NLW_$1I4585/NC_O_UNCONNECTED ;
  wire \NLW_$1I4586/NC_O_UNCONNECTED ;
  wire \NLW_$1I4587/NC_O_UNCONNECTED ;
  wire \NLW_$1I4588/NC_O_UNCONNECTED ;
  wire \NLW_$1I4589/NC_O_UNCONNECTED ;
  wire \NLW_$1I4590/NC_O_UNCONNECTED ;
  wire \NLW_$1I4591/NC_O_UNCONNECTED ;
  wire \NLW_$1I4592/NC_O_UNCONNECTED ;
  wire \NLW_$1I4593/NC_O_UNCONNECTED ;
  wire \NLW_$1I4594/NC_O_UNCONNECTED ;
  wire \NLW_$1I4595/NC_O_UNCONNECTED ;
  wire \NLW_$1I4596/NC_O_UNCONNECTED ;
  wire \NLW_$1I4597/NC_O_UNCONNECTED ;
  wire \NLW_$1I4598/NC_O_UNCONNECTED ;
  wire \NLW_$1I4599/NC_O_UNCONNECTED ;
  wire \NLW_$1I4600/NC_O_UNCONNECTED ;
  wire \NLW_$1I4601/NC_O_UNCONNECTED ;
  wire \NLW_$1I4602/NC_O_UNCONNECTED ;
  wire \NLW_$1I4603/NC_O_UNCONNECTED ;
  wire \NLW_$1I4604/NC_O_UNCONNECTED ;
  wire \NLW_$1I4605/NC_O_UNCONNECTED ;
  wire \NLW_$1I4606/NC_O_UNCONNECTED ;
  wire \NLW_$1I4607/NC_O_UNCONNECTED ;
  wire \NLW_$1I4608/NC_O_UNCONNECTED ;
  wire \NLW_$1I4609/NC_O_UNCONNECTED ;
  wire \NLW_$1I4610/NC_O_UNCONNECTED ;
  wire \NlwInverterSignal_TDLY/$1I315/M01/$1I31/I0 ;
  wire \NlwInverterSignal_TDLY/$1I315/M23/$1I31/I0 ;
  wire \NlwInverterSignal_TDLY/$1I328/M01/$1I31/I0 ;
  wire \NlwInverterSignal_TDLY/$1I328/M23/$1I31/I0 ;
  wire \NlwInverterSignal_IDLY/$1I315/M01/$1I31/I0 ;
  wire \NlwInverterSignal_IDLY/$1I315/M23/$1I31/I0 ;
  wire \NlwInverterSignal_IDLY/$1I328/M01/$1I31/I0 ;
  wire \NlwInverterSignal_IDLY/$1I328/M23/$1I31/I0 ;
  wire \NlwInverterSignal_DATA_VLD/$1I426/I0 ;
  wire \NlwInverterSignal_DATA_VLD/$1I426/I1 ;
  wire \NlwInverterSignal_DATA_VLD/$1I328/I0 ;
  wire \NlwInverterSignal_DATA_VLD/$1I328/I1 ;
  wire \NlwInverterSignal_SRC_EN/$1I742/I0 ;
  wire \NlwInverterSignal_SRC_EN/$1I656/I0 ;
  wire \NlwInverterSignal_SRC_EN/$1I615/I0 ;
  wire \NlwInverterSignal_SRC_EN/$1I558/I0 ;
  wire \NLW_SRC_EN/$1I736/NC_O_UNCONNECTED ;
  wire \NLW_SRC_EN/$1I737/NC_O_UNCONNECTED ;
  wire \NlwInverterSignal_OUT_CE/$3I1079/I0 ;
  wire \NlwInverterSignal_OUT_CE/$3I1079/O ;
  wire \NlwInverterSignal_OUT_CE/$3I1078/I0 ;
  wire \NlwInverterSignal_OUT_CE/$3I1078/O ;
  wire \NlwInverterSignal_OUT_CE/$3I1062/I0 ;
  wire \NlwInverterSignal_OUT_CE/$3I1062/I1 ;
  wire \NlwInverterSignal_OUT_CE/$3I1061/I0 ;
  wire \NlwInverterSignal_OUT_CE/$3I1061/I1 ;
  wire \NlwInverterSignal_OUT_CE/$3I1056/I0 ;
  wire \NlwInverterSignal_OUT_CE/$2I1086/I0 ;
  wire \NlwInverterSignal_OUT_CE/$2I1086/I1 ;
  wire \NlwInverterSignal_OUT_CE/$2I1085/I0 ;
  wire \NlwInverterSignal_OUT_CE/$2I1085/I1 ;
  wire \NlwInverterSignal_OUT_CE/$2I1084/I0 ;
  wire \NlwInverterSignal_OUT_CE/$2I1084/I1 ;
  wire \NlwInverterSignal_OUT_CE/$2I1083/I0 ;
  wire \NlwInverterSignal_OUT_CE/$2I1083/I1 ;
  wire \NlwInverterSignal_OUT_CE/$2I1015/I0 ;
  wire \NlwInverterSignal_OUT_CE/$2I1015/I1 ;
  wire \NlwInverterSignal_OUT_CE/$2I1013/I0 ;
  wire \NlwInverterSignal_OUT_CE/$2I1013/I1 ;
  wire \NlwInverterSignal_OUT_CE/$2I1012/I0 ;
  wire \NlwInverterSignal_OUT_CE/$2I1012/I1 ;
  wire \NlwInverterSignal_OUT_CE/$2I1007/I0 ;
  wire \NlwInverterSignal_OUT_CE/$2I1007/I1 ;
  wire \NlwInverterSignal_OUT_CE/$1I980/I0 ;
  wire \NlwInverterSignal_OUT_CE/$1I976/I0 ;
  wire \NlwInverterSignal_OUT_CE/$1I975/I0 ;
  wire \NlwInverterSignal_OUT_CE/$1I972/I0 ;
  wire \NlwInverterSignal_OUT_CE/MAGICBOX/PCI_CE/I0 ;
  wire \NlwInverterSignal_OUT_CE/MAGICBOX/PCI_CE/O ;
  wire \NlwInverterSignal_OUT_CE/MAGICBOX/I3_NAND_TRDY/I0 ;
  wire \NlwInverterSignal_OUT_CE/MAGICBOX/I3_NAND_TRDY/I1 ;
  wire \NlwInverterSignal_OUT_CE/MAGICBOX/I3_NAND_TRDY/O ;
  wire \NlwInverterSignal_OUT_CE/MAGICBOX/I1_NAND_IRDY/I0 ;
  wire \NlwInverterSignal_OUT_CE/MAGICBOX/I1_NAND_IRDY/I1 ;
  wire \NlwInverterSignal_OUT_CE/MAGICBOX/I1_NAND_IRDY/O ;
  wire \NlwInverterSignal_OUT_CE/$4I1005/$1I7/I0 ;
  wire \NlwInverterSignal_OUT_SEL/$1I916/I0 ;
  wire \NlwInverterSignal_OUT_SEL/$1I916/I1 ;
  wire \NlwInverterSignal_OUT_SEL/$1I913/I0 ;
  wire \NlwInverterSignal_OUT_SEL/$1I913/I1 ;
  wire \NlwInverterSignal_OUT_SEL/$1I913/I2 ;
  wire \NlwInverterSignal_OUT_SEL/$1I897/I0 ;
  wire \NlwInverterSignal_OUT_SEL/$1I853/I0 ;
  wire \NlwInverterSignal_OUT_SEL/$1I849/I0 ;
  wire \NlwInverterSignal_OUT_SEL/$1I758/I0 ;
  wire \NlwInverterSignal_ADDR_VLD/$1I4008/I0 ;
  wire \NlwInverterSignal_ADDR_VLD/$1I4008/I1 ;
  wire \NlwInverterSignal_ADDR_VLD/$1I4005/I0 ;
  wire \NlwInverterSignal_ADDR_VLD/$1I4005/O ;
  wire \NlwInverterSignal_ADDR_VLD/$1I3989/I0 ;
  wire \NlwInverterSignal_ADDR_VLD/$1I3989/O ;
  wire \NlwInverterSignal_ADDR_VLD/$1I3986/I0 ;
  wire \NlwInverterSignal_ADDR_VLD/$1I3986/O ;
  wire \NlwInverterSignal_ADDR_VLD/$1I3983/I0 ;
  wire \NlwInverterSignal_ADDR_VLD/$1I3983/O ;
  wire \NlwInverterSignal_ADDR_VLD/$1I3980/I0 ;
  wire \NlwInverterSignal_ADDR_VLD/$1I3980/O ;
  wire \NlwInverterSignal_ADDR_VLD/$1I3963/I0 ;
  wire \NlwInverterSignal_ADDR_VLD/$1I3894/I0 ;
  wire \NlwInverterSignal_ADDR_VLD/$1I3880/I0 ;
  wire \NlwInverterSignal_ADDR_VLD/$1I3867/I0 ;
  wire \NlwInverterSignal_EOT/$1I617/I0 ;
  wire \NlwInverterSignal_EOT/$1I617/I1 ;
  wire \NlwInverterSignal_EOT/$1I616/I0 ;
  wire \NlwInverterSignal_EOT/$1I615/I0 ;
  wire \NlwInverterSignal_EOT/$1I615/I1 ;
  wire \NlwInverterSignal_EOT/$1I589/I0 ;
  wire \NlwInverterSignal_EOT/$1I589/I1 ;
  wire \NlwInverterSignal_EOT/$1I588/I0 ;
  wire \NlwInverterSignal_PCI-PAR/$7I2985/O ;
  wire \NlwInverterSignal_PCI-PAR/$7I2974/O ;
  wire \NlwInverterSignal_PCI-PAR/$4I3127/O ;
  wire \NlwInverterSignal_PCI-PAR/$4I3104/O ;
  wire \NlwInverterSignal_PCI-PAR/$3I3057/I0 ;
  wire \NlwInverterSignal_PCI-PAR/$3I3018/O ;
  wire \NlwInverterSignal_PCI-PAR/$3I2993/O ;
  wire \NlwInverterSignal_PCI-PAR/$3I2940/O ;
  wire \NlwInverterSignal_PCI-PAR/$3I2936/I0 ;
  wire \NlwInverterSignal_PCI-PAR/$3I2931/I0 ;
  wire \NlwInverterSignal_4/UPPER/T0/T ;
  wire \NlwInverterSignal_4/UPPER/T1/T ;
  wire \NlwInverterSignal_4/UPPER/T2/T ;
  wire \NlwInverterSignal_4/UPPER/T3/T ;
  wire \NlwInverterSignal_4/UPPER/T4/T ;
  wire \NlwInverterSignal_4/UPPER/T5/T ;
  wire \NlwInverterSignal_4/UPPER/T6/T ;
  wire \NlwInverterSignal_4/UPPER/T7/T ;
  wire \NlwInverterSignal_4/UPPER/T8/T ;
  wire \NlwInverterSignal_4/UPPER/T9/T ;
  wire \NlwInverterSignal_4/UPPER/T10/T ;
  wire \NlwInverterSignal_4/UPPER/T11/T ;
  wire \NlwInverterSignal_4/UPPER/T12/T ;
  wire \NlwInverterSignal_4/UPPER/T13/T ;
  wire \NlwInverterSignal_4/UPPER/T14/T ;
  wire \NlwInverterSignal_4/UPPER/T15/T ;
  wire \NlwInverterSignal_4/LOWER/T0/T ;
  wire \NlwInverterSignal_4/LOWER/T1/T ;
  wire \NlwInverterSignal_4/LOWER/T2/T ;
  wire \NlwInverterSignal_4/LOWER/T3/T ;
  wire \NlwInverterSignal_4/LOWER/T4/T ;
  wire \NlwInverterSignal_4/LOWER/T5/T ;
  wire \NlwInverterSignal_4/LOWER/T6/T ;
  wire \NlwInverterSignal_4/LOWER/T7/T ;
  wire \NlwInverterSignal_4/LOWER/T8/T ;
  wire \NlwInverterSignal_4/LOWER/T9/T ;
  wire \NlwInverterSignal_4/LOWER/T10/T ;
  wire \NlwInverterSignal_4/LOWER/T11/T ;
  wire \NlwInverterSignal_4/LOWER/T12/T ;
  wire \NlwInverterSignal_4/LOWER/T13/T ;
  wire \NlwInverterSignal_4/LOWER/T14/T ;
  wire \NlwInverterSignal_4/LOWER/T15/T ;
  wire \NlwInverterSignal_5/UPPER/T0/T ;
  wire \NlwInverterSignal_5/UPPER/T1/T ;
  wire \NlwInverterSignal_5/UPPER/T2/T ;
  wire \NlwInverterSignal_5/UPPER/T3/T ;
  wire \NlwInverterSignal_5/UPPER/T4/T ;
  wire \NlwInverterSignal_5/UPPER/T5/T ;
  wire \NlwInverterSignal_5/UPPER/T6/T ;
  wire \NlwInverterSignal_5/UPPER/T7/T ;
  wire \NlwInverterSignal_5/UPPER/T8/T ;
  wire \NlwInverterSignal_5/UPPER/T9/T ;
  wire \NlwInverterSignal_5/UPPER/T10/T ;
  wire \NlwInverterSignal_5/UPPER/T11/T ;
  wire \NlwInverterSignal_5/UPPER/T12/T ;
  wire \NlwInverterSignal_5/UPPER/T13/T ;
  wire \NlwInverterSignal_5/UPPER/T14/T ;
  wire \NlwInverterSignal_5/UPPER/T15/T ;
  wire \NlwInverterSignal_5/LOWER/T0/T ;
  wire \NlwInverterSignal_5/LOWER/T1/T ;
  wire \NlwInverterSignal_5/LOWER/T2/T ;
  wire \NlwInverterSignal_5/LOWER/T3/T ;
  wire \NlwInverterSignal_5/LOWER/T4/T ;
  wire \NlwInverterSignal_5/LOWER/T5/T ;
  wire \NlwInverterSignal_5/LOWER/T6/T ;
  wire \NlwInverterSignal_5/LOWER/T7/T ;
  wire \NlwInverterSignal_5/LOWER/T8/T ;
  wire \NlwInverterSignal_5/LOWER/T9/T ;
  wire \NlwInverterSignal_5/LOWER/T10/T ;
  wire \NlwInverterSignal_5/LOWER/T11/T ;
  wire \NlwInverterSignal_5/LOWER/T12/T ;
  wire \NlwInverterSignal_5/LOWER/T13/T ;
  wire \NlwInverterSignal_5/LOWER/T14/T ;
  wire \NlwInverterSignal_5/LOWER/T15/T ;
  wire \NlwInverterSignal_6/UPPER/T0/T ;
  wire \NlwInverterSignal_6/UPPER/T1/T ;
  wire \NlwInverterSignal_6/UPPER/T2/T ;
  wire \NlwInverterSignal_6/UPPER/T3/T ;
  wire \NlwInverterSignal_6/UPPER/T4/T ;
  wire \NlwInverterSignal_6/UPPER/T5/T ;
  wire \NlwInverterSignal_6/UPPER/T6/T ;
  wire \NlwInverterSignal_6/UPPER/T7/T ;
  wire \NlwInverterSignal_6/UPPER/T8/T ;
  wire \NlwInverterSignal_6/UPPER/T9/T ;
  wire \NlwInverterSignal_6/UPPER/T10/T ;
  wire \NlwInverterSignal_6/UPPER/T11/T ;
  wire \NlwInverterSignal_6/UPPER/T12/T ;
  wire \NlwInverterSignal_6/UPPER/T13/T ;
  wire \NlwInverterSignal_6/UPPER/T14/T ;
  wire \NlwInverterSignal_6/UPPER/T15/T ;
  wire \NlwInverterSignal_6/LOWER/T0/T ;
  wire \NlwInverterSignal_6/LOWER/T1/T ;
  wire \NlwInverterSignal_6/LOWER/T2/T ;
  wire \NlwInverterSignal_6/LOWER/T3/T ;
  wire \NlwInverterSignal_6/LOWER/T4/T ;
  wire \NlwInverterSignal_6/LOWER/T5/T ;
  wire \NlwInverterSignal_6/LOWER/T6/T ;
  wire \NlwInverterSignal_6/LOWER/T7/T ;
  wire \NlwInverterSignal_6/LOWER/T8/T ;
  wire \NlwInverterSignal_6/LOWER/T9/T ;
  wire \NlwInverterSignal_6/LOWER/T10/T ;
  wire \NlwInverterSignal_6/LOWER/T11/T ;
  wire \NlwInverterSignal_6/LOWER/T12/T ;
  wire \NlwInverterSignal_6/LOWER/T13/T ;
  wire \NlwInverterSignal_6/LOWER/T14/T ;
  wire \NlwInverterSignal_6/LOWER/T15/T ;
  wire \NLW_$3I3818/NC_O_UNCONNECTED ;
  wire \NLW_$3I3819/NC_O_UNCONNECTED ;
  wire \NLW_$3I3820/NC_O_UNCONNECTED ;
  wire \NLW_$3I3821/NC_O_UNCONNECTED ;
  wire \NLW_$3I3822/NC_O_UNCONNECTED ;
  wire \NLW_$3I3823/NC_O_UNCONNECTED ;
  wire \NLW_$3I3824/NC_O_UNCONNECTED ;
  wire \NLW_$3I3825/NC_O_UNCONNECTED ;
  wire \NLW_$3I3826/NC_O_UNCONNECTED ;
  wire \NLW_$3I3827/NC_O_UNCONNECTED ;
  wire \NLW_$3I3828/NC_O_UNCONNECTED ;
  wire \NLW_$3I3829/NC_O_UNCONNECTED ;
  wire \NLW_$3I3830/NC_O_UNCONNECTED ;
  wire \NLW_$3I3831/NC_O_UNCONNECTED ;
  wire \NLW_$3I3832/NC_O_UNCONNECTED ;
  wire \NLW_$3I3833/NC_O_UNCONNECTED ;
  wire \NlwInverterSignal_BAR0/BR-31-24/X1/O ;
  wire \NlwInverterSignal_BAR0/BR-31-24/X3/O ;
  wire \NlwInverterSignal_BAR0/BR-31-24/X2/O ;
  wire \NlwInverterSignal_BAR0/BR-31-24/X0/O ;
  wire \NlwInverterSignal_BAR0/BR-31-24/X4/O ;
  wire \NlwInverterSignal_BAR0/BR-31-24/X6/O ;
  wire \NlwInverterSignal_BAR0/BR-31-24/X7/O ;
  wire \NlwInverterSignal_BAR0/BR-31-24/X5/O ;
  wire \NlwInverterSignal_BAR0/BR-23-16/X1/O ;
  wire \NlwInverterSignal_BAR0/BR-23-16/X3/O ;
  wire \NlwInverterSignal_BAR0/BR-23-16/X2/O ;
  wire \NlwInverterSignal_BAR0/BR-23-16/X0/O ;
  wire \NlwInverterSignal_BAR0/BR-23-16/X4/O ;
  wire \NlwInverterSignal_BAR0/BR-23-16/X6/O ;
  wire \NlwInverterSignal_BAR0/BR-23-16/X7/O ;
  wire \NlwInverterSignal_BAR0/BR-23-16/X5/O ;
  wire \NlwInverterSignal_BAR0/BR-15-8/X1/O ;
  wire \NlwInverterSignal_BAR0/BR-15-8/X3/O ;
  wire \NlwInverterSignal_BAR0/BR-15-8/X2/O ;
  wire \NlwInverterSignal_BAR0/BR-15-8/X0/O ;
  wire \NlwInverterSignal_BAR0/BR-15-8/X4/O ;
  wire \NlwInverterSignal_BAR0/BR-15-8/X6/O ;
  wire \NlwInverterSignal_BAR0/BR-15-8/X7/O ;
  wire \NlwInverterSignal_BAR0/BR-15-8/X5/O ;
  wire \NlwInverterSignal_BAR0/BR-CMD/$1I194/I0 ;
  wire \NlwInverterSignal_BAR0/BR-CMD/$1I173/I0 ;
  wire \NlwInverterSignal_BAR0/BR-CMD/$1I173/I1 ;
  wire \NlwInverterSignal_BAR0/BR-CMD/$1I117/I0 ;
  wire \NlwInverterSignal_BAR0/BR-CMD/$1I110/I0 ;
  wire \NlwInverterSignal_BAR0/BR-CMD/$1I100/I0 ;
  wire \NlwInverterSignal_BAR0/BR-CMD/$1I223/$1I31/I0 ;
  wire \NlwInverterSignal_BAR0/BR-7-4/X7/O ;
  wire \NlwInverterSignal_BAR0/BR-7-4/X6/O ;
  wire \NlwInverterSignal_BAR0/BR-7-4/X5/O ;
  wire \NlwInverterSignal_BAR0/BR-7-4/X4/O ;
  wire \NlwInverterSignal_BAR0/$1I3440/$1I31/I0 ;
  wire \NlwInverterSignal_BAR0/$1I3453/$1I31/I0 ;
  wire \NlwInverterSignal_BAR0/$2I3321/$1I31/I0 ;
  wire \NlwInverterSignal_BAR1/BR-31-24/X1/O ;
  wire \NlwInverterSignal_BAR1/BR-31-24/X3/O ;
  wire \NlwInverterSignal_BAR1/BR-31-24/X2/O ;
  wire \NlwInverterSignal_BAR1/BR-31-24/X0/O ;
  wire \NlwInverterSignal_BAR1/BR-31-24/X4/O ;
  wire \NlwInverterSignal_BAR1/BR-31-24/X6/O ;
  wire \NlwInverterSignal_BAR1/BR-31-24/X7/O ;
  wire \NlwInverterSignal_BAR1/BR-31-24/X5/O ;
  wire \NlwInverterSignal_BAR1/BR-23-16/X1/O ;
  wire \NlwInverterSignal_BAR1/BR-23-16/X3/O ;
  wire \NlwInverterSignal_BAR1/BR-23-16/X2/O ;
  wire \NlwInverterSignal_BAR1/BR-23-16/X0/O ;
  wire \NlwInverterSignal_BAR1/BR-23-16/X4/O ;
  wire \NlwInverterSignal_BAR1/BR-23-16/X6/O ;
  wire \NlwInverterSignal_BAR1/BR-23-16/X7/O ;
  wire \NlwInverterSignal_BAR1/BR-23-16/X5/O ;
  wire \NlwInverterSignal_BAR1/BR-15-8/X1/O ;
  wire \NlwInverterSignal_BAR1/BR-15-8/X3/O ;
  wire \NlwInverterSignal_BAR1/BR-15-8/X2/O ;
  wire \NlwInverterSignal_BAR1/BR-15-8/X0/O ;
  wire \NlwInverterSignal_BAR1/BR-15-8/X4/O ;
  wire \NlwInverterSignal_BAR1/BR-15-8/X6/O ;
  wire \NlwInverterSignal_BAR1/BR-15-8/X7/O ;
  wire \NlwInverterSignal_BAR1/BR-15-8/X5/O ;
  wire \NlwInverterSignal_BAR1/BR-CMD/$1I194/I0 ;
  wire \NlwInverterSignal_BAR1/BR-CMD/$1I173/I0 ;
  wire \NlwInverterSignal_BAR1/BR-CMD/$1I173/I1 ;
  wire \NlwInverterSignal_BAR1/BR-CMD/$1I117/I0 ;
  wire \NlwInverterSignal_BAR1/BR-CMD/$1I110/I0 ;
  wire \NlwInverterSignal_BAR1/BR-CMD/$1I100/I0 ;
  wire \NlwInverterSignal_BAR1/BR-CMD/$1I223/$1I31/I0 ;
  wire \NlwInverterSignal_BAR1/BR-7-4/X7/O ;
  wire \NlwInverterSignal_BAR1/BR-7-4/X6/O ;
  wire \NlwInverterSignal_BAR1/BR-7-4/X5/O ;
  wire \NlwInverterSignal_BAR1/BR-7-4/X4/O ;
  wire \NlwInverterSignal_BAR1/$1I3440/$1I31/I0 ;
  wire \NlwInverterSignal_BAR1/$1I3453/$1I31/I0 ;
  wire \NlwInverterSignal_BAR1/$2I3321/$1I31/I0 ;
  wire \NlwInverterSignal_BAR2/BR-31-24/X1/O ;
  wire \NlwInverterSignal_BAR2/BR-31-24/X3/O ;
  wire \NlwInverterSignal_BAR2/BR-31-24/X2/O ;
  wire \NlwInverterSignal_BAR2/BR-31-24/X0/O ;
  wire \NlwInverterSignal_BAR2/BR-31-24/X4/O ;
  wire \NlwInverterSignal_BAR2/BR-31-24/X6/O ;
  wire \NlwInverterSignal_BAR2/BR-31-24/X7/O ;
  wire \NlwInverterSignal_BAR2/BR-31-24/X5/O ;
  wire \NlwInverterSignal_BAR2/BR-23-16/X1/O ;
  wire \NlwInverterSignal_BAR2/BR-23-16/X3/O ;
  wire \NlwInverterSignal_BAR2/BR-23-16/X2/O ;
  wire \NlwInverterSignal_BAR2/BR-23-16/X0/O ;
  wire \NlwInverterSignal_BAR2/BR-23-16/X4/O ;
  wire \NlwInverterSignal_BAR2/BR-23-16/X6/O ;
  wire \NlwInverterSignal_BAR2/BR-23-16/X7/O ;
  wire \NlwInverterSignal_BAR2/BR-23-16/X5/O ;
  wire \NlwInverterSignal_BAR2/BR-15-8/X1/O ;
  wire \NlwInverterSignal_BAR2/BR-15-8/X3/O ;
  wire \NlwInverterSignal_BAR2/BR-15-8/X2/O ;
  wire \NlwInverterSignal_BAR2/BR-15-8/X0/O ;
  wire \NlwInverterSignal_BAR2/BR-15-8/X4/O ;
  wire \NlwInverterSignal_BAR2/BR-15-8/X6/O ;
  wire \NlwInverterSignal_BAR2/BR-15-8/X7/O ;
  wire \NlwInverterSignal_BAR2/BR-15-8/X5/O ;
  wire \NlwInverterSignal_BAR2/BR-CMD/$1I194/I0 ;
  wire \NlwInverterSignal_BAR2/BR-CMD/$1I173/I0 ;
  wire \NlwInverterSignal_BAR2/BR-CMD/$1I173/I1 ;
  wire \NlwInverterSignal_BAR2/BR-CMD/$1I117/I0 ;
  wire \NlwInverterSignal_BAR2/BR-CMD/$1I110/I0 ;
  wire \NlwInverterSignal_BAR2/BR-CMD/$1I100/I0 ;
  wire \NlwInverterSignal_BAR2/BR-CMD/$1I223/$1I31/I0 ;
  wire \NlwInverterSignal_BAR2/BR-7-4/X7/O ;
  wire \NlwInverterSignal_BAR2/BR-7-4/X6/O ;
  wire \NlwInverterSignal_BAR2/BR-7-4/X5/O ;
  wire \NlwInverterSignal_BAR2/BR-7-4/X4/O ;
  wire \NlwInverterSignal_BAR2/$1I3440/$1I31/I0 ;
  wire \NlwInverterSignal_BAR2/$1I3453/$1I31/I0 ;
  wire \NlwInverterSignal_BAR2/$2I3321/$1I31/I0 ;
  wire \NlwInverterSignal_F/UPPER/T0/T ;
  wire \NlwInverterSignal_F/UPPER/T1/T ;
  wire \NlwInverterSignal_F/UPPER/T2/T ;
  wire \NlwInverterSignal_F/UPPER/T3/T ;
  wire \NlwInverterSignal_F/UPPER/T4/T ;
  wire \NlwInverterSignal_F/UPPER/T5/T ;
  wire \NlwInverterSignal_F/UPPER/T6/T ;
  wire \NlwInverterSignal_F/UPPER/T7/T ;
  wire \NlwInverterSignal_F/UPPER/T8/T ;
  wire \NlwInverterSignal_F/UPPER/T9/T ;
  wire \NlwInverterSignal_F/UPPER/T10/T ;
  wire \NlwInverterSignal_F/UPPER/T11/T ;
  wire \NlwInverterSignal_F/UPPER/T12/T ;
  wire \NlwInverterSignal_F/UPPER/T13/T ;
  wire \NlwInverterSignal_F/UPPER/T14/T ;
  wire \NlwInverterSignal_F/UPPER/T15/T ;
  wire \NlwInverterSignal_F/LOWER/T0/T ;
  wire \NlwInverterSignal_F/LOWER/T1/T ;
  wire \NlwInverterSignal_F/LOWER/T2/T ;
  wire \NlwInverterSignal_F/LOWER/T3/T ;
  wire \NlwInverterSignal_F/LOWER/T4/T ;
  wire \NlwInverterSignal_F/LOWER/T5/T ;
  wire \NlwInverterSignal_F/LOWER/T6/T ;
  wire \NlwInverterSignal_F/LOWER/T7/T ;
  wire \NlwInverterSignal_F/LOWER/T8/T ;
  wire \NlwInverterSignal_F/LOWER/T9/T ;
  wire \NlwInverterSignal_F/LOWER/T10/T ;
  wire \NlwInverterSignal_F/LOWER/T11/T ;
  wire \NlwInverterSignal_F/LOWER/T12/T ;
  wire \NlwInverterSignal_F/LOWER/T13/T ;
  wire \NlwInverterSignal_F/LOWER/T14/T ;
  wire \NlwInverterSignal_F/LOWER/T15/T ;
  wire \NlwInverterSignal_1/UPPER/T0/T ;
  wire \NlwInverterSignal_1/UPPER/T1/T ;
  wire \NlwInverterSignal_1/UPPER/T2/T ;
  wire \NlwInverterSignal_1/UPPER/T3/T ;
  wire \NlwInverterSignal_1/UPPER/T4/T ;
  wire \NlwInverterSignal_1/UPPER/T5/T ;
  wire \NlwInverterSignal_1/UPPER/T6/T ;
  wire \NlwInverterSignal_1/UPPER/T7/T ;
  wire \NlwInverterSignal_1/UPPER/T8/T ;
  wire \NlwInverterSignal_1/UPPER/T9/T ;
  wire \NlwInverterSignal_1/UPPER/T10/T ;
  wire \NlwInverterSignal_1/UPPER/T11/T ;
  wire \NlwInverterSignal_1/UPPER/T12/T ;
  wire \NlwInverterSignal_1/UPPER/T13/T ;
  wire \NlwInverterSignal_1/UPPER/T14/T ;
  wire \NlwInverterSignal_1/UPPER/T15/T ;
  wire \NlwInverterSignal_1/LOWER/T0/T ;
  wire \NlwInverterSignal_1/LOWER/T1/T ;
  wire \NlwInverterSignal_1/LOWER/T2/T ;
  wire \NlwInverterSignal_1/LOWER/T3/T ;
  wire \NlwInverterSignal_1/LOWER/T4/T ;
  wire \NlwInverterSignal_1/LOWER/T5/T ;
  wire \NlwInverterSignal_1/LOWER/T6/T ;
  wire \NlwInverterSignal_1/LOWER/T7/T ;
  wire \NlwInverterSignal_1/LOWER/T8/T ;
  wire \NlwInverterSignal_1/LOWER/T9/T ;
  wire \NlwInverterSignal_1/LOWER/T10/T ;
  wire \NlwInverterSignal_1/LOWER/T11/T ;
  wire \NlwInverterSignal_1/LOWER/T12/T ;
  wire \NlwInverterSignal_1/LOWER/T13/T ;
  wire \NlwInverterSignal_1/LOWER/T14/T ;
  wire \NlwInverterSignal_1/LOWER/T15/T ;
  wire \NlwInverterSignal_0/UPPER/T0/T ;
  wire \NlwInverterSignal_0/UPPER/T1/T ;
  wire \NlwInverterSignal_0/UPPER/T2/T ;
  wire \NlwInverterSignal_0/UPPER/T3/T ;
  wire \NlwInverterSignal_0/UPPER/T4/T ;
  wire \NlwInverterSignal_0/UPPER/T5/T ;
  wire \NlwInverterSignal_0/UPPER/T6/T ;
  wire \NlwInverterSignal_0/UPPER/T7/T ;
  wire \NlwInverterSignal_0/UPPER/T8/T ;
  wire \NlwInverterSignal_0/UPPER/T9/T ;
  wire \NlwInverterSignal_0/UPPER/T10/T ;
  wire \NlwInverterSignal_0/UPPER/T11/T ;
  wire \NlwInverterSignal_0/UPPER/T12/T ;
  wire \NlwInverterSignal_0/UPPER/T13/T ;
  wire \NlwInverterSignal_0/UPPER/T14/T ;
  wire \NlwInverterSignal_0/UPPER/T15/T ;
  wire \NlwInverterSignal_0/LOWER/T0/T ;
  wire \NlwInverterSignal_0/LOWER/T1/T ;
  wire \NlwInverterSignal_0/LOWER/T2/T ;
  wire \NlwInverterSignal_0/LOWER/T3/T ;
  wire \NlwInverterSignal_0/LOWER/T4/T ;
  wire \NlwInverterSignal_0/LOWER/T5/T ;
  wire \NlwInverterSignal_0/LOWER/T6/T ;
  wire \NlwInverterSignal_0/LOWER/T7/T ;
  wire \NlwInverterSignal_0/LOWER/T8/T ;
  wire \NlwInverterSignal_0/LOWER/T9/T ;
  wire \NlwInverterSignal_0/LOWER/T10/T ;
  wire \NlwInverterSignal_0/LOWER/T11/T ;
  wire \NlwInverterSignal_0/LOWER/T12/T ;
  wire \NlwInverterSignal_0/LOWER/T13/T ;
  wire \NlwInverterSignal_0/LOWER/T14/T ;
  wire \NlwInverterSignal_0/LOWER/T15/T ;
  wire \NLW_PCI-IREG/$1I2521/NC_O_UNCONNECTED ;
  wire \NLW_PCI-IREG/$1I2555/NC_O_UNCONNECTED ;
  wire \NLW_PCI-IREG/$1I2557/NC_O_UNCONNECTED ;
  wire \NLW_PCI-IREG/$1I2559/NC_O_UNCONNECTED ;
  wire \NLW_PCI-IREG/$1I2561/NC_O_UNCONNECTED ;
  wire \NLW_PCI-IREG/$1I2563/NC_O_UNCONNECTED ;
  wire \NLW_PCI-IREG/$1I2565/NC_O_UNCONNECTED ;
  wire \NLW_PCI-IREG/$1I2567/NC_O_UNCONNECTED ;
  wire \NLW_PCI-IREG/$1I2569/NC_O_UNCONNECTED ;
  wire \NLW_PCI-IREG/$1I2582/NC_O_UNCONNECTED ;
  wire \NLW_PCI-IREG/$1I2584/NC_O_UNCONNECTED ;
  wire \NLW_PCI-CSR/CMDREG/$1I2492/NC_O_UNCONNECTED ;
  wire \NLW_PCI-CSR/CMDREG/$1I2495/NC_O_UNCONNECTED ;
  wire \NLW_PCI-CSR/CMDREG/$1I2497/NC_O_UNCONNECTED ;
  wire \NLW_PCI-CSR/CMDREG/$1I2499/NC_O_UNCONNECTED ;
  wire \NLW_PCI-CSR/CMDREG/$1I2501/NC_O_UNCONNECTED ;
  wire \NLW_PCI-CSR/CMDREG/$1I2505/NC_O_UNCONNECTED ;
  wire \NLW_PCI-CSR/CMDREG/$1I2507/NC_O_UNCONNECTED ;
  wire \NLW_PCI-CSR/CMDREG/$1I2509/NC_O_UNCONNECTED ;
  wire \NLW_PCI-CSR/CMDREG/$1I2538/NC_O_UNCONNECTED ;
  wire \NLW_PCI-CSR/CMDREG/$1I2540/NC_O_UNCONNECTED ;
  wire \NLW_PCI-CSR/CMDREG/$1I2551/NC_O_UNCONNECTED ;
  wire \NLW_PCI-CSR/CMDREG/$1I2552/NC_O_UNCONNECTED ;
  wire \NlwInverterSignal_PCI-CSR/STATREG/Q14/$1I2230/I0 ;
  wire \NlwInverterSignal_PCI-CSR/STATREG/Q14/$1I2233/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-CSR/STATREG/Q12/$1I2230/I0 ;
  wire \NlwInverterSignal_PCI-CSR/STATREG/Q12/$1I2233/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-CSR/STATREG/Q8/$1I2230/I0 ;
  wire \NlwInverterSignal_PCI-CSR/STATREG/Q8/$1I2233/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-CSR/STATREG/Q11/$1I2230/I0 ;
  wire \NlwInverterSignal_PCI-CSR/STATREG/Q11/$1I2233/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-CSR/STATREG/Q13/$1I2230/I0 ;
  wire \NlwInverterSignal_PCI-CSR/STATREG/Q13/$1I2233/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-CSR/STATREG/Q15/$1I2230/I0 ;
  wire \NlwInverterSignal_PCI-CSR/STATREG/Q15/$1I2233/$1I7/I0 ;
  wire \NLW_PCI-CSR/STATREG/$1I2497/NC_O_UNCONNECTED ;
  wire \NLW_PCI-CSR/STATREG/$1I2500/NC_O_UNCONNECTED ;
  wire \NLW_PCI-CSR/STATREG/$1I2502/NC_O_UNCONNECTED ;
  wire \NLW_PCI-CSR/STATREG/$1I2504/NC_O_UNCONNECTED ;
  wire \NLW_PCI-CSR/STATREG/$1I2506/NC_O_UNCONNECTED ;
  wire \NLW_PCI-CSR/STATREG/$1I2508/NC_O_UNCONNECTED ;
  wire \NLW_PCI-CSR/STATREG/$1I2510/NC_O_UNCONNECTED ;
  wire \NLW_PCI-CSR/STATREG/$1I2512/NC_O_UNCONNECTED ;
  wire \NLW_PCI-CSR/STATREG/$1I2514/NC_O_UNCONNECTED ;
  wire \NLW_PCI-CSR/STATREG/$1I2523/NC_O_UNCONNECTED ;
  wire \NLW_PCI-CSR/STATREG/$1I2524/NC_O_UNCONNECTED ;
  wire \NLW_PCI-CSR/STATREG/$1I2525/NC_O_UNCONNECTED ;
  wire \NLW_PCI-CSR/STATREG/$1I2526/NC_O_UNCONNECTED ;
  wire \NLW_PCI-CSR/STATREG/$1I2527/NC_O_UNCONNECTED ;
  wire \NLW_PCI-CSR/STATREG/$1I2528/NC_O_UNCONNECTED ;
  wire \NLW_PCI-CSR/STATREG/$1I2529/NC_O_UNCONNECTED ;
  wire \NLW_PCI-CSR/STATREG/$1I2530/NC_O_UNCONNECTED ;
  wire \NLW_PCI-CSR/STATREG/$1I2532/NC_O_UNCONNECTED ;
  wire \NLW_PCI-CSR/STATREG/$1I2598/NC_O_UNCONNECTED ;
  wire \NLW_PCI-CSR/STATREG/$1I2600/NC_O_UNCONNECTED ;
  wire \NLW_PCI-CSR/STATREG/$1I2612/NC_O_UNCONNECTED ;
  wire \NLW_PCI-CSR/STATREG/$1I2613/NC_O_UNCONNECTED ;
  wire \NlwInverterSignal_PCI-ROM/$1I8330/I0 ;
  wire \NlwInverterSignal_PCI-ROM/$1I8330/I1 ;
  wire \NlwInverterSignal_PCI-ROM/$1I8282/I0 ;
  wire \NlwInverterSignal_PCI-ROM/$1I8282/I1 ;
  wire \NlwInverterSignal_PCI-ROM/$1I8282/I2 ;
  wire \NlwInverterSignal_PCI-ROM/$1I8237/I0 ;
  wire \NlwInverterSignal_PCI-ROM/$1I8237/I1 ;
  wire \NlwInverterSignal_PCI-ROM/$1I8227/I0 ;
  wire \NlwInverterSignal_PCI-ROM/$1I8227/I1 ;
  wire \NlwInverterSignal_PCI-ROM/$1I8227/I2 ;
  wire \NlwInverterSignal_PCI-ROM/$1I8110/I0 ;
  wire \NlwInverterSignal_PCI-ROM/$1I8110/I1 ;
  wire \NlwInverterSignal_PCI-ROM/$1I8078/I0 ;
  wire \NlwInverterSignal_PCI-ROM/$1I8078/I1 ;
  wire \NLW_PCI-ROM/$1I8479/NC_O_UNCONNECTED ;
  wire \NLW_PCI-ROM/$1I8480/NC_O_UNCONNECTED ;
  wire \NLW_PCI-ROM/$1I8481/NC_O_UNCONNECTED ;
  wire \NLW_PCI-ROM/$1I8482/NC_O_UNCONNECTED ;
  wire \NLW_PCI-ROM/$1I8483/NC_O_UNCONNECTED ;
  wire \NLW_PCI-ROM/$1I8484/NC_O_UNCONNECTED ;
  wire \NLW_PCI-ROM/$1I8485/NC_O_UNCONNECTED ;
  wire \NLW_PCI-ROM/$1I8486/NC_O_UNCONNECTED ;
  wire \NLW_PCI-ROM/$1I8487/NC_O_UNCONNECTED ;
  wire \NLW_PCI-ROM/$1I8488/NC_O_UNCONNECTED ;
  wire \NLW_PCI-ROM/$1I8489/NC_O_UNCONNECTED ;
  wire \NLW_PCI-ROM/$1I8490/NC_O_UNCONNECTED ;
  wire \NLW_PCI-ROM/$1I8491/NC_O_UNCONNECTED ;
  wire \NLW_PCI-ROM/$1I8492/NC_O_UNCONNECTED ;
  wire \NLW_PCI-ROM/$1I8493/NC_O_UNCONNECTED ;
  wire \NLW_PCI-ROM/$1I8494/NC_O_UNCONNECTED ;
  wire \NLW_PCI-ROM/$1I8495/NC_O_UNCONNECTED ;
  wire \NLW_PCI-ROM/$1I8496/NC_O_UNCONNECTED ;
  wire \NLW_PCI-ROM/$1I8497/NC_O_UNCONNECTED ;
  wire \NLW_PCI-ROM/$1I8498/NC_O_UNCONNECTED ;
  wire \NLW_PCI-ROM/$1I8499/NC_O_UNCONNECTED ;
  wire \NLW_PCI-ROM/$1I8500/NC_O_UNCONNECTED ;
  wire \NLW_PCI-ROM/$1I8501/NC_O_UNCONNECTED ;
  wire \NLW_PCI-ROM/$1I8502/NC_O_UNCONNECTED ;
  wire \NLW_PCI-ROM/$1I8503/NC_O_UNCONNECTED ;
  wire \NLW_PCI-ROM/$1I8504/NC_O_UNCONNECTED ;
  wire \NLW_PCI-ROM/$1I8505/NC_O_UNCONNECTED ;
  wire \NLW_PCI-ROM/$1I8506/NC_O_UNCONNECTED ;
  wire \NLW_PCI-ROM/$1I8507/NC_O_UNCONNECTED ;
  wire \NLW_PCI-ROM/$1I8508/NC_O_UNCONNECTED ;
  wire \NLW_PCI-ROM/$1I8509/NC_O_UNCONNECTED ;
  wire \NLW_PCI-ROM/$1I8510/NC_O_UNCONNECTED ;
  wire \NlwInverterSignal_$4I4029/$1I2610/$1I43/$1I30/$1I7/I0 ;
  wire \NlwInverterSignal_$4I4029/$1I2610/$1I53/$1I30/$1I7/I0 ;
  wire \NlwInverterSignal_$4I4029/$1I2610/$1I58/$1I30/$1I7/I0 ;
  wire \NlwInverterSignal_$4I4029/$1I2610/$1I59/$1I30/$1I7/I0 ;
  wire \NlwInverterSignal_$4I4029/$1I2610/$1I68/$1I30/$1I7/I0 ;
  wire \NlwInverterSignal_$4I4029/$1I2610/$1I73/$1I30/$1I7/I0 ;
  wire \NlwInverterSignal_$4I4029/$1I2610/$1I79/$1I30/$1I7/I0 ;
  wire \NlwInverterSignal_$4I4029/$1I2610/$1I84/$1I30/$1I7/I0 ;
  wire \NlwInverterSignal_$4I4029/$1I2637/$1I43/$1I30/$1I7/I0 ;
  wire \NlwInverterSignal_$4I4029/$1I2637/$1I53/$1I30/$1I7/I0 ;
  wire \NlwInverterSignal_$4I4029/$1I2637/$1I58/$1I30/$1I7/I0 ;
  wire \NlwInverterSignal_$4I4029/$1I2637/$1I59/$1I30/$1I7/I0 ;
  wire \NlwInverterSignal_$4I4029/$1I2637/$1I68/$1I30/$1I7/I0 ;
  wire \NlwInverterSignal_$4I4029/$1I2637/$1I73/$1I30/$1I7/I0 ;
  wire \NlwInverterSignal_$4I4029/$1I2637/$1I79/$1I30/$1I7/I0 ;
  wire \NlwInverterSignal_$4I4029/$1I2637/$1I84/$1I30/$1I7/I0 ;
  wire \NlwInverterSignal_$4I4029/$1I2645/$1I43/$1I30/$1I7/I0 ;
  wire \NlwInverterSignal_$4I4029/$1I2645/$1I53/$1I30/$1I7/I0 ;
  wire \NlwInverterSignal_$4I4029/$1I2645/$1I58/$1I30/$1I7/I0 ;
  wire \NlwInverterSignal_$4I4029/$1I2645/$1I59/$1I30/$1I7/I0 ;
  wire \NlwInverterSignal_$4I4029/$1I2645/$1I68/$1I30/$1I7/I0 ;
  wire \NlwInverterSignal_$4I4029/$1I2645/$1I73/$1I30/$1I7/I0 ;
  wire \NlwInverterSignal_$4I4029/$1I2645/$1I79/$1I30/$1I7/I0 ;
  wire \NlwInverterSignal_$4I4029/$1I2645/$1I84/$1I30/$1I7/I0 ;
  wire \NlwInverterSignal_$4I4029/$1I2653/$1I43/$1I30/$1I7/I0 ;
  wire \NlwInverterSignal_$4I4029/$1I2653/$1I53/$1I30/$1I7/I0 ;
  wire \NlwInverterSignal_$4I4029/$1I2653/$1I58/$1I30/$1I7/I0 ;
  wire \NlwInverterSignal_$4I4029/$1I2653/$1I59/$1I30/$1I7/I0 ;
  wire \NlwInverterSignal_$4I4029/$1I2653/$1I68/$1I30/$1I7/I0 ;
  wire \NlwInverterSignal_$4I4029/$1I2653/$1I73/$1I30/$1I7/I0 ;
  wire \NlwInverterSignal_$4I4029/$1I2653/$1I79/$1I30/$1I7/I0 ;
  wire \NlwInverterSignal_$4I4029/$1I2653/$1I84/$1I30/$1I7/I0 ;
  wire \NlwInverterSignal_$4I4029/$1I2661/$1I43/$1I30/$1I7/I0 ;
  wire \NlwInverterSignal_$4I4029/$1I2661/$1I53/$1I30/$1I7/I0 ;
  wire \NlwInverterSignal_$4I4029/$1I2661/$1I58/$1I30/$1I7/I0 ;
  wire \NlwInverterSignal_$4I4029/$1I2661/$1I59/$1I30/$1I7/I0 ;
  wire \NlwInverterSignal_$4I4029/$1I2661/$1I68/$1I30/$1I7/I0 ;
  wire \NlwInverterSignal_$4I4029/$1I2661/$1I73/$1I30/$1I7/I0 ;
  wire \NlwInverterSignal_$4I4029/$1I2661/$1I79/$1I30/$1I7/I0 ;
  wire \NlwInverterSignal_$4I4029/$1I2661/$1I84/$1I30/$1I7/I0 ;
  wire \NlwInverterSignal_E/UPPER/T0/T ;
  wire \NlwInverterSignal_E/UPPER/T1/T ;
  wire \NlwInverterSignal_E/UPPER/T2/T ;
  wire \NlwInverterSignal_E/UPPER/T3/T ;
  wire \NlwInverterSignal_E/UPPER/T4/T ;
  wire \NlwInverterSignal_E/UPPER/T5/T ;
  wire \NlwInverterSignal_E/UPPER/T6/T ;
  wire \NlwInverterSignal_E/UPPER/T7/T ;
  wire \NlwInverterSignal_E/UPPER/T8/T ;
  wire \NlwInverterSignal_E/UPPER/T9/T ;
  wire \NlwInverterSignal_E/UPPER/T10/T ;
  wire \NlwInverterSignal_E/UPPER/T11/T ;
  wire \NlwInverterSignal_E/UPPER/T12/T ;
  wire \NlwInverterSignal_E/UPPER/T13/T ;
  wire \NlwInverterSignal_E/UPPER/T14/T ;
  wire \NlwInverterSignal_E/UPPER/T15/T ;
  wire \NlwInverterSignal_E/LOWER/T0/T ;
  wire \NlwInverterSignal_E/LOWER/T1/T ;
  wire \NlwInverterSignal_E/LOWER/T2/T ;
  wire \NlwInverterSignal_E/LOWER/T3/T ;
  wire \NlwInverterSignal_E/LOWER/T4/T ;
  wire \NlwInverterSignal_E/LOWER/T5/T ;
  wire \NlwInverterSignal_E/LOWER/T6/T ;
  wire \NlwInverterSignal_E/LOWER/T7/T ;
  wire \NlwInverterSignal_E/LOWER/T8/T ;
  wire \NlwInverterSignal_E/LOWER/T9/T ;
  wire \NlwInverterSignal_E/LOWER/T10/T ;
  wire \NlwInverterSignal_E/LOWER/T11/T ;
  wire \NlwInverterSignal_E/LOWER/T12/T ;
  wire \NlwInverterSignal_E/LOWER/T13/T ;
  wire \NlwInverterSignal_E/LOWER/T14/T ;
  wire \NlwInverterSignal_E/LOWER/T15/T ;
  wire \NlwInverterSignal_E64/UPPER/T0/T ;
  wire \NlwInverterSignal_E64/UPPER/T1/T ;
  wire \NlwInverterSignal_E64/UPPER/T2/T ;
  wire \NlwInverterSignal_E64/UPPER/T3/T ;
  wire \NlwInverterSignal_E64/UPPER/T4/T ;
  wire \NlwInverterSignal_E64/UPPER/T5/T ;
  wire \NlwInverterSignal_E64/UPPER/T6/T ;
  wire \NlwInverterSignal_E64/UPPER/T7/T ;
  wire \NlwInverterSignal_E64/UPPER/T8/T ;
  wire \NlwInverterSignal_E64/UPPER/T9/T ;
  wire \NlwInverterSignal_E64/UPPER/T10/T ;
  wire \NlwInverterSignal_E64/UPPER/T11/T ;
  wire \NlwInverterSignal_E64/UPPER/T12/T ;
  wire \NlwInverterSignal_E64/UPPER/T13/T ;
  wire \NlwInverterSignal_E64/UPPER/T14/T ;
  wire \NlwInverterSignal_E64/UPPER/T15/T ;
  wire \NlwInverterSignal_E64/LOWER/T0/T ;
  wire \NlwInverterSignal_E64/LOWER/T1/T ;
  wire \NlwInverterSignal_E64/LOWER/T2/T ;
  wire \NlwInverterSignal_E64/LOWER/T3/T ;
  wire \NlwInverterSignal_E64/LOWER/T4/T ;
  wire \NlwInverterSignal_E64/LOWER/T5/T ;
  wire \NlwInverterSignal_E64/LOWER/T6/T ;
  wire \NlwInverterSignal_E64/LOWER/T7/T ;
  wire \NlwInverterSignal_E64/LOWER/T8/T ;
  wire \NlwInverterSignal_E64/LOWER/T9/T ;
  wire \NlwInverterSignal_E64/LOWER/T10/T ;
  wire \NlwInverterSignal_E64/LOWER/T11/T ;
  wire \NlwInverterSignal_E64/LOWER/T12/T ;
  wire \NlwInverterSignal_E64/LOWER/T13/T ;
  wire \NlwInverterSignal_E64/LOWER/T14/T ;
  wire \NlwInverterSignal_E64/LOWER/T15/T ;
  wire \NlwInverterSignal_OEADI/$1I4041/I0 ;
  wire \NlwInverterSignal_OEADI/$1I4040/I0 ;
  wire \NlwInverterSignal_OEADI/$1I4031/I0 ;
  wire \NlwInverterSignal_OEADI/$1I4031/I1 ;
  wire \NlwInverterSignal_OEADI/$1I4031/I2 ;
  wire \NlwInverterSignal_OEADI/$1I4031/O ;
  wire \NlwInverterSignal_OEADI/$1I4028/I0 ;
  wire \NlwInverterSignal_OEADI/$1I4028/O ;
  wire \NlwInverterSignal_OEADI/$1I3984/I0 ;
  wire \NlwInverterSignal_OEADI/$1I3984/O ;
  wire \NlwInverterSignal_OEADI/$1I3954/I0 ;
  wire \NlwInverterSignal_OEADI/$1I3954/I1 ;
  wire \NlwInverterSignal_OEADI/$1I3954/I2 ;
  wire \NlwInverterSignal_OEADI/$1I3954/O ;
  wire \NlwInverterSignal_OEADI/$1I3864/I0 ;
  wire \NlwInverterSignal_OEADI/$1I3860/I0 ;
  wire \NLW_OEADI/$1I4047/NC_O_UNCONNECTED ;
  wire \NlwInverterSignal_$5I3771/$1I7/I0 ;
  wire \NlwInverterSignal_$5I3781/$1I7/I0 ;
  wire \NLW_$6I1087/NC_O_UNCONNECTED ;
  wire \NLW_$6I1090/NC_O_UNCONNECTED ;
  wire \NlwInverterSignal_DEVSEL/$1I2310/M01/$1I31/I0 ;
  wire \NlwInverterSignal_DEVSEL/$1I2310/M23/$1I31/I0 ;
  wire \NlwInverterSignal_ACK64/$1I2310/M01/$1I31/I0 ;
  wire \NlwInverterSignal_ACK64/$1I2310/M23/$1I31/I0 ;
  wire \NlwInverterSignal_FRAME/$1I2310/M01/$1I31/I0 ;
  wire \NlwInverterSignal_FRAME/$1I2310/M23/$1I31/I0 ;
  wire \NlwInverterSignal_TRDY/$1I2310/M01/$1I31/I0 ;
  wire \NlwInverterSignal_TRDY/$1I2310/M23/$1I31/I0 ;
  wire \NlwInverterSignal_REQ64/$1I2310/M01/$1I31/I0 ;
  wire \NlwInverterSignal_REQ64/$1I2310/M23/$1I31/I0 ;
  wire \NlwInverterSignal_IRDY/$1I2310/M01/$1I31/I0 ;
  wire \NlwInverterSignal_IRDY/$1I2310/M23/$1I31/I0 ;
  wire \NlwInverterSignal_STOP/$1I2310/M01/$1I31/I0 ;
  wire \NlwInverterSignal_STOP/$1I2310/M23/$1I31/I0 ;
  wire \NlwInverterSignal_$7I576/$1I7/I0 ;
  wire \NlwInverterSignal_$7I577/$1I7/I0 ;
  wire \NlwInverterSignal_$7I622/$1I7/I0 ;
  wire \NlwInverterSignal_$7I623/$1I7/I0 ;
  wire \NlwInverterSignal_$7I824/$1I7/I0 ;
  wire \NlwInverterSignal_$7I826/$1I7/I0 ;
  wire \NlwInverterSignal_$7I828/$1I7/I0 ;
  wire \NlwInverterSignal_$7I830/$1I7/I0 ;
  wire \NlwInverterSignal_$7I832/$1I7/I0 ;
  wire \NlwInverterSignal_$7I834/$1I7/I0 ;
  wire \NlwInverterSignal_$7I836/$1I7/I0 ;
  wire \NlwInverterSignal_$7I838/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-CBE/$1I2773/I0 ;
  wire \NlwInverterSignal_PCI-CBE/IO3/$1I2296/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-CBE/IO3/$1I2303/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-CBE/IO2/$1I2296/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-CBE/IO2/$1I2303/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-CBE/IO1/$1I2296/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-CBE/IO1/$1I2303/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-CBE/IO0/$1I2296/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-CBE/IO0/$1I2303/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-CBE/$1I2777/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-CBE/$1I2779/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/IO28/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/IO30/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/IO29/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/IO31/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/IO20/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/IO22/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/IO21/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/IO23/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/IO12/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/IO14/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/IO13/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/IO15/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/IO4/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/IO6/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/IO5/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/IO7/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/$1I2927/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/$1I2928/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/$1I2929/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/$1I2930/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/$1I2931/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/$1I2932/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/$1I2933/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/$1I2934/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/$1I2935/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/$1I2936/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/$1I2937/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/$1I2938/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/$1I2939/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/$1I2940/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/$1I2941/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/$1I2942/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/$1I2943/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/$1I2944/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/$1I2945/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/$1I2946/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/$1I2947/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/$1I2948/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/$1I2949/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/$1I2950/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/$1I2951/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/$1I2952/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/$1I2953/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/$1I2954/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/$1I2955/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/$1I2956/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/$1I2957/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/$1I2958/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/IO27/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/IO26/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/IO25/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/IO24/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/IO19/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/IO18/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/IO17/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/IO16/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/IO11/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/IO10/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/IO9/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/IO8/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/IO3/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/IO2/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/IO1/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD/IO0/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD64/IO28/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD64/IO30/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD64/IO29/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD64/IO31/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD64/IO20/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD64/IO22/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD64/IO21/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD64/IO23/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD64/IO12/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD64/IO14/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD64/IO13/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD64/IO15/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD64/IO4/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD64/IO6/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD64/IO5/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD64/IO7/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD64/IO27/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD64/IO26/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD64/IO25/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD64/IO24/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD64/IO19/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD64/IO18/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD64/IO17/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD64/IO16/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD64/IO11/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD64/IO10/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD64/IO9/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD64/IO8/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD64/IO3/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD64/IO2/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD64/IO1/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-AD64/IO0/$1I2246/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-CBE64/IO3/$1I2296/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-CBE64/IO3/$1I2303/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-CBE64/IO2/$1I2296/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-CBE64/IO2/$1I2303/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-CBE64/IO1/$1I2296/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-CBE64/IO1/$1I2303/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-CBE64/IO0/$1I2296/$1I7/I0 ;
  wire \NlwInverterSignal_PCI-CBE64/IO0/$1I2303/$1I7/I0 ;
  assign
    BASE_HIT0 = NlwRenamedSig_OI_BASE_HIT0,
    BASE_HIT1 = NlwRenamedSig_OI_BASE_HIT1,
    BASE_HIT2 = NlwRenamedSig_OI_BASE_HIT2,
    BASE_HIT3 = NlwRenamedSig_OI_BASE_HIT3,
    BASE_HIT4 = NlwRenamedSig_OI_BASE_HIT4,
    BASE_HIT5 = NlwRenamedSig_OI_BASE_HIT5,
    BASE_HIT6 = NlwRenamedSig_OI_BASE_HIT6,
    BASE_HIT7 = NlwRenamedSig_OI_BASE_HIT7,
    OE_CBE = NlwRenamedSig_OI_OE_CBE,
    OE_ADO_LT64 = NlwRenamedSig_OI_OE_ADO_LT64,
    CSR10 = NlwRenamedSig_OI_CSR10,
    CSR11 = NlwRenamedSig_OI_CSR11,
    CSR12 = NlwRenamedSig_OI_CSR12,
    CSR13 = NlwRenamedSig_OI_CSR13,
    CSR14 = NlwRenamedSig_OI_CSR14,
    CSR15 = NlwRenamedSig_OI_CSR15,
    CSR16 = NlwRenamedSig_OI_CSR16,
    CSR20 = NlwRenamedSig_OI_CSR20,
    CSR17 = NlwRenamedSig_OI_CSR17,
    CSR21 = NlwRenamedSig_OI_CSR21,
    CSR18 = NlwRenamedSig_OI_CSR18,
    CSR22 = NlwRenamedSig_OI_CSR22,
    CSR19 = NlwRenamedSig_OI_CSR19,
    CSR23 = NlwRenamedSig_OI_CSR23,
    CSR24 = NlwRenamedSig_OI_CSR24,
    CSR25 = NlwRenamedSig_OI_CSR25,
    CSR26 = NlwRenamedSig_OI_CSR26,
    CSR30 = NlwRenamedSig_OI_CSR30,
    CSR27 = NlwRenamedSig_OI_CSR27,
    CSR31 = NlwRenamedSig_OI_CSR31,
    CSR28 = NlwRenamedSig_OI_CSR28,
    CSR32 = NlwRenamedSig_OI_CSR32,
    CSR29 = NlwRenamedSig_OI_CSR29,
    CSR33 = NlwRenamedSig_OI_CSR33,
    CSR34 = NlwRenamedSig_OI_CSR34,
    CSR35 = NlwRenamedSig_OI_CSR35,
    CSR36 = NlwRenamedSig_OI_CSR36,
    CSR37 = NlwRenamedSig_OI_CSR37,
    CSR38 = NlwRenamedSig_OI_CSR38,
    CSR39 = NlwRenamedSig_OI_CSR39,
    PCI_CMD0 = NlwRenamedSig_OI_PCI_CMD0,
    PCI_CMD1 = NlwRenamedSig_OI_PCI_CMD1,
    PCI_CMD2 = NlwRenamedSig_OI_PCI_CMD2,
    PCI_CMD3 = NlwRenamedSig_OI_PCI_CMD3,
    PCI_CMD4 = NlwRenamedSig_OI_PCI_CMD4,
    PCI_CMD5 = NlwRenamedSig_OI_PCI_CMD5,
    PCI_CMD6 = NlwRenamedSig_OI_PCI_CMD6,
    PCI_CMD7 = NlwRenamedSig_OI_PCI_CMD7,
    PCI_CMD8 = NlwRenamedSig_OI_PCI_CMD8,
    PCI_CMD9 = NlwRenamedSig_OI_PCI_CMD9,
    S_CBE0 = NlwRenamedSig_OI_S_CBE0,
    S_CBE1 = NlwRenamedSig_OI_S_CBE1,
    S_CBE2 = NlwRenamedSig_OI_S_CBE2,
    S_CBE3 = NlwRenamedSig_OI_S_CBE3,
    ADDR_VLD = NlwRenamedSig_OI_ADDR_VLD,
    S_CBE4 = NlwRenamedSig_OI_S_CBE4,
    S_CBE5 = NlwRenamedSig_OI_S_CBE5,
    S_CBE6 = NlwRenamedSig_OI_S_CBE6,
    S_CBE7 = NlwRenamedSig_OI_S_CBE7,
    S_WRDN = NlwRenamedSig_OI_S_WRDN,
    RST = NlwRenamedSig_OI_RST,
    PCI_CMD10 = NlwRenamedSig_OI_PCI_CMD10,
    PCI_CMD11 = NlwRenamedSig_OI_PCI_CMD11,
    PCI_CMD12 = NlwRenamedSig_OI_PCI_CMD12,
    PCI_CMD13 = NlwRenamedSig_OI_PCI_CMD13,
    PCI_CMD14 = NlwRenamedSig_OI_PCI_CMD14,
    PCI_CMD15 = NlwRenamedSig_OI_PCI_CMD15,
    CSR0 = NlwRenamedSig_OI_CSR0,
    CSR1 = NlwRenamedSig_OI_CSR1,
    CSR2 = NlwRenamedSig_OI_CSR2,
    CSR3 = NlwRenamedSig_OI_CSR3,
    CSR4 = NlwRenamedSig_OI_CSR4,
    CSR5 = NlwRenamedSig_OI_CSR5,
    CSR6 = NlwRenamedSig_OI_CSR6,
    CSR7 = NlwRenamedSig_OI_CSR7,
    CSR8 = NlwRenamedSig_OI_CSR8,
    CSR9 = NlwRenamedSig_OI_CSR9,
    ADDR10 = NlwRenamedSig_OI_ADDR10,
    ADDR11 = NlwRenamedSig_OI_ADDR11,
    ADDR12 = NlwRenamedSig_OI_ADDR12,
    ADDR13 = NlwRenamedSig_OI_ADDR13,
    ADDR14 = NlwRenamedSig_OI_ADDR14,
    ADDR15 = NlwRenamedSig_OI_ADDR15,
    ADDR16 = NlwRenamedSig_OI_ADDR16,
    ADDR20 = NlwRenamedSig_OI_ADDR20,
    ADDR17 = NlwRenamedSig_OI_ADDR17,
    ADDR21 = NlwRenamedSig_OI_ADDR21,
    ADDR18 = NlwRenamedSig_OI_ADDR18,
    ADDR22 = NlwRenamedSig_OI_ADDR22,
    ADDR19 = NlwRenamedSig_OI_ADDR19,
    ADDR23 = NlwRenamedSig_OI_ADDR23,
    ADDR24 = NlwRenamedSig_OI_ADDR24,
    ADDR25 = NlwRenamedSig_OI_ADDR25,
    ADDR26 = NlwRenamedSig_OI_ADDR26,
    ADDR30 = NlwRenamedSig_OI_ADDR30,
    ADDR27 = NlwRenamedSig_OI_ADDR27,
    ADDR31 = NlwRenamedSig_OI_ADDR31,
    ADDR28 = NlwRenamedSig_OI_ADDR28,
    ADDR29 = NlwRenamedSig_OI_ADDR29,
    OE_ADO_B = NlwRenamedSig_OI_OE_ADO_B,
    M_SRC_EN = NlwRenamedSig_OI_M_SRC_EN,
    OE_ADO_T = NlwRenamedSig_OI_OE_ADO_T,
    TIME_OUT = NlwRenamedSig_OI_TIME_OUT,
    OE_ADO_B64 = NlwRenamedSig_OI_OE_ADO_B64,
    CFG_VLD = NlwRenamedSig_OI_CFG_VLD,
    OE_PAR = NlwRenamedSig_OI_OE_PAR,
    OE_ADO_LB64 = NlwRenamedSig_OI_OE_ADO_LB64,
    ADDR0 = NlwRenamedSig_OI_ADDR0,
    OE_PAR64 = NlwRenamedSig_OI_OE_PAR64,
    ADDR1 = NlwRenamedSig_OI_ADDR1,
    ADDR2 = NlwRenamedSig_OI_ADDR2,
    ADDR3 = NlwRenamedSig_OI_ADDR3,
    ADDR4 = NlwRenamedSig_OI_ADDR4,
    ADDR5 = NlwRenamedSig_OI_ADDR5,
    ADDR6 = NlwRenamedSig_OI_ADDR6,
    ADDR7 = NlwRenamedSig_OI_ADDR7,
    ADDR8 = NlwRenamedSig_OI_ADDR8,
    OE_ADO_T64 = NlwRenamedSig_OI_OE_ADO_T64,
    ADDR9 = NlwRenamedSig_OI_ADDR9,
    CFG_HIT = NlwRenamedSig_OI_CFG_HIT,
    OE_CBE64 = NlwRenamedSig_OI_OE_CBE64,
    OE_ADO_LB = NlwRenamedSig_OI_OE_ADO_LB,
    OE_ADO_LT = NlwRenamedSig_OI_OE_ADO_LT;
  X_INV   \$1I4832  (
    .I(CFG249),
    .O(\$1N4834 )
  );
  X_BUF   \$3I3130  (
    .I(BAR7),
    .O(NlwRenamedSig_OI_BASE_HIT7)
  );
  X_BUF   \$3I3131  (
    .I(BAR6),
    .O(NlwRenamedSig_OI_BASE_HIT6)
  );
  X_BUF   \$3I3132  (
    .I(BAR5),
    .O(NlwRenamedSig_OI_BASE_HIT5)
  );
  X_BUF   \$3I3133  (
    .I(BAR4),
    .O(NlwRenamedSig_OI_BASE_HIT4)
  );
  X_BUF   \$3I3134  (
    .I(BAR3),
    .O(NlwRenamedSig_OI_BASE_HIT3)
  );
  X_BUF   \$3I3349  (
    .I(NL7),
    .O(NL_MEM7)
  );
  X_BUF   \$3I3350  (
    .I(NL6),
    .O(NL_MEM6)
  );
  X_BUF   \$3I3351  (
    .I(NL5),
    .O(NL_MEM5)
  );
  X_BUF   \$3I3352  (
    .I(NL4),
    .O(NL_MEM4)
  );
  X_BUF   \$3I3353  (
    .I(NL3),
    .O(NL_MEM3)
  );
  X_OR2   \$3I3487  (
    .I0(\NlwInverterSignal_$3I3487/I0 ),
    .I1(OE4),
    .O(BAR0_T)
  );
  X_OR2   \$3I3492  (
    .I0(\NlwInverterSignal_$3I3492/I0 ),
    .I1(OE5),
    .O(BAR1_T)
  );
  X_OR2   \$3I3496  (
    .I0(\NlwInverterSignal_$3I3496/I0 ),
    .I1(OE6),
    .O(BAR2_T)
  );
  X_AND2   \$4I4017  (
    .I0(\NlwInverterSignal_$4I4017/I0 ),
    .I1(\NlwInverterSignal_$4I4017/I1 ),
    .O(\NlwInverterSignal_$4I4017/O )
  );
  X_OR2   \$5I3767  (
    .I0(CFG252),
    .I1(OE_ADI64),
    .O(DP64_T)
  );
  X_INV   \$6I1083  (
    .I(RST_N),
    .O(NlwRenamedSig_OI_RST)
  );
  X_AND2   \$6I1164  (
    .I0(CFG73),
    .I1(CFG37),
    .O(\$6N1152 )
  );
  X_AND2   \$6I1165  (
    .I0(CFG36),
    .I1(CFG0),
    .O(\$6N1151 )
  );
  X_OR3   \$6I1166  (
    .I0(\$6N1153 ),
    .I1(\$6N1152 ),
    .I2(\$6N1151 ),
    .O(HAS_IO)
  );
  X_OR3   \$6I1167  (
    .I0(\$6N1154 ),
    .I1(\$6N1155 ),
    .I2(\$6N1156 ),
    .O(HAS_MEM)
  );
  X_AND3   \$6I1168  (
    .I0(\NlwInverterSignal_$6I1168/I0 ),
    .I1(\NlwInverterSignal_$6I1168/I1 ),
    .I2(CFG74),
    .O(\$6N1154 )
  );
  X_AND2   \$6I1169  (
    .I0(\NlwInverterSignal_$6I1169/I0 ),
    .I1(CFG37),
    .O(\$6N1155 )
  );
  X_AND3   \$6I1170  (
    .I0(\NlwInverterSignal_$6I1170/I0 ),
    .I1(CFG110),
    .I2(CFG74),
    .O(\$6N1153 )
  );
  X_AND2   \$6I1172  (
    .I0(\NlwInverterSignal_$6I1172/I0 ),
    .I1(CFG0),
    .O(\$6N1156 )
  );
  X_AND2   \$7I129  (
    .I0(\NlwInverterSignal_$7I129/I0 ),
    .I1(\NlwInverterSignal_$7I129/I1 ),
    .O(\$7N147 )
  );
  X_AND3   \$7I130  (
    .I0(\NlwInverterSignal_$7I130/I0 ),
    .I1(\FRAME- ),
    .I2(\STOP- ),
    .O(\$7N149 )
  );
  X_AND2   \$7I131  (
    .I0(\NlwInverterSignal_$7I131/I0 ),
    .I1(\FRAME- ),
    .O(\$7N152 )
  );
  X_AND3   \$7I132  (
    .I0(\NlwInverterSignal_$7I132/I0 ),
    .I1(\NlwInverterSignal_$7I132/I1 ),
    .I2(\TRDY- ),
    .O(\$7N156 )
  );
  X_AND3   \$7I133  (
    .I0(\NlwInverterSignal_$7I133/I0 ),
    .I1(\NlwInverterSignal_$7I133/I1 ),
    .I2(\NlwInverterSignal_$7I133/I2 ),
    .O(\$7N160 )
  );
  X_AND2   \$7I134  (
    .I0(\NlwInverterSignal_$7I134/I0 ),
    .I1(\DEVSEL- ),
    .O(\$7N163 )
  );
  X_AND2   \$7I140  (
    .I0(\$7N143 ),
    .I1(\FRAME- ),
    .O(\$7N148 )
  );
  X_OR2   \$7I141  (
    .I0(\NlwInverterSignal_$7I141/I0 ),
    .I1(\NlwInverterSignal_$7I141/I1 ),
    .O(\$7N143 )
  );
  X_BUF   \$7I427  (
    .I(\FRAME- ),
    .O(FRAMEQ_N)
  );
  X_BUF   \$7I431  (
    .I(\IRDY- ),
    .O(IRDYQ_N)
  );
  X_BUF   \$7I434  (
    .I(\DEVSEL- ),
    .O(DEVSELQ_N)
  );
  X_BUF   \$7I437  (
    .I(\TRDY- ),
    .O(TRDYQ_N)
  );
  X_BUF   \$7I440  (
    .I(\STOP- ),
    .O(STOPQ_N)
  );
  X_BUF   \$7I476  (
    .I(\PERR- ),
    .O(PERRQ_N)
  );
  X_BUF   \$7I490  (
    .I(S_CYCLE64_INT),
    .O(S_CYCLE64)
  );
  X_BUF   \$7I493  (
    .I(IDLE_INT),
    .O(IDLE)
  );
  X_BUF   \$7I496  (
    .I(B_BUSY_INT),
    .O(B_BUSY)
  );
  X_BUF   \$7I502  (
    .I(I_IDLE_INT),
    .O(I_IDLE)
  );
  X_BUF   \$7I505  (
    .I(DR_BUS_INT),
    .O(DR_BUS)
  );
  X_BUF   \$7I600  (
    .I(\REQ64- ),
    .O(REQ64Q_N)
  );
  X_BUF   \$7I618  (
    .I(\ACK64- ),
    .O(ACK64Q_N)
  );
  X_BUF   \$7I701  (
    .I(NlwRenamedSig_OI_CSR2),
    .O(M_ENABLE)
  );
  X_BUF   \$7I702  (
    .I(NlwRenamedSig_OI_CSR6),
    .O(PERR_EN)
  );
  X_BUF   \$7I703  (
    .I(NlwRenamedSig_OI_CSR8),
    .O(SERR_EN)
  );
  X_BUF   \$7I724  (
    .I(CBE_IN7),
    .O(NlwRenamedSig_OI_S_CBE7)
  );
  X_BUF   \$7I725  (
    .I(CBE_IN6),
    .O(NlwRenamedSig_OI_S_CBE6)
  );
  X_BUF   \$7I726  (
    .I(CBE_IN5),
    .O(NlwRenamedSig_OI_S_CBE5)
  );
  X_BUF   \$7I727  (
    .I(CBE_IN4),
    .O(NlwRenamedSig_OI_S_CBE4)
  );
  X_BUF   \$7I728  (
    .I(CBE_IN3),
    .O(NlwRenamedSig_OI_S_CBE3)
  );
  X_BUF   \$7I729  (
    .I(CBE_IN2),
    .O(NlwRenamedSig_OI_S_CBE2)
  );
  X_BUF   \$7I730  (
    .I(CBE_IN1),
    .O(NlwRenamedSig_OI_S_CBE1)
  );
  X_BUF   \$7I731  (
    .I(CBE_IN0),
    .O(NlwRenamedSig_OI_S_CBE0)
  );
  X_BUF   \$7I734  (
    .I(\SERR- ),
    .O(SERRQ_N)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \$7I737  (
    .CE(VCC),
    .CLK(CLK),
    .I(INTACK),
    .O(INTACKQ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b1 ))
  FAKE_GTS (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(CLK),
    .I(\$7N745 ),
    .O(FAKE_GTS_13003),
    .RST(GND)
  );
  X_BUF   \$7I753  (
    .I(FAIL64_INT),
    .O(M_FAIL64)
  );
  X_OR2   \$7I792  (
    .I0(FAKE_GTS_13003),
    .I1(M_CBE7),
    .O(M_CBE_INT7)
  );
  X_OR2   \$7I793  (
    .I0(FAKE_GTS_13003),
    .I1(M_CBE6),
    .O(M_CBE_INT6)
  );
  X_OR2   \$7I794  (
    .I0(FAKE_GTS_13003),
    .I1(M_CBE5),
    .O(M_CBE_INT5)
  );
  X_OR2   \$7I795  (
    .I0(FAKE_GTS_13003),
    .I1(M_CBE4),
    .O(M_CBE_INT4)
  );
  X_OR2   \$7I796  (
    .I0(FAKE_GTS_13003),
    .I1(M_CBE3),
    .O(M_CBE_INT3)
  );
  X_OR2   \$7I797  (
    .I0(FAKE_GTS_13003),
    .I1(M_CBE2),
    .O(M_CBE_INT2)
  );
  X_OR2   \$7I798  (
    .I0(FAKE_GTS_13003),
    .I1(M_CBE1),
    .O(M_CBE_INT1)
  );
  X_OR2   \$7I799  (
    .I0(FAKE_GTS_13003),
    .I1(M_CBE0),
    .O(M_CBE_INT0)
  );
  X_BUF   \$7I806  (
    .I(BACKOFF_INT),
    .O(BACKOFF)
  );
  X_AND3   \$7I863  (
    .I0(\NlwInverterSignal_$7I863/I0 ),
    .I1(NlwRenamedSig_OI_ADDR_VLD),
    .I2(\$7N583 ),
    .O(INTACK)
  );
  X_PU   \ADIO0.PULLUP  (
    .O(ADIO0)
  );
  X_PU   \ADIO1.PULLUP  (
    .O(ADIO1)
  );
  X_PU   \ADIO10.PULLUP  (
    .O(ADIO10)
  );
  X_PU   \ADIO11.PULLUP  (
    .O(ADIO11)
  );
  X_PU   \ADIO12.PULLUP  (
    .O(ADIO12)
  );
  X_PU   \ADIO13.PULLUP  (
    .O(ADIO13)
  );
  X_PU   \ADIO14.PULLUP  (
    .O(ADIO14)
  );
  X_PU   \ADIO15.PULLUP  (
    .O(ADIO15)
  );
  X_PU   \ADIO16.PULLUP  (
    .O(ADIO16)
  );
  X_PU   \ADIO17.PULLUP  (
    .O(ADIO17)
  );
  X_PU   \ADIO18.PULLUP  (
    .O(ADIO18)
  );
  X_PU   \ADIO19.PULLUP  (
    .O(ADIO19)
  );
  X_PU   \ADIO2.PULLUP  (
    .O(ADIO2)
  );
  X_PU   \ADIO20.PULLUP  (
    .O(ADIO20)
  );
  X_PU   \ADIO21.PULLUP  (
    .O(ADIO21)
  );
  X_PU   \ADIO22.PULLUP  (
    .O(ADIO22)
  );
  X_PU   \ADIO23.PULLUP  (
    .O(ADIO23)
  );
  X_PU   \ADIO24.PULLUP  (
    .O(ADIO24)
  );
  X_PU   \ADIO25.PULLUP  (
    .O(ADIO25)
  );
  X_PU   \ADIO26.PULLUP  (
    .O(ADIO26)
  );
  X_PU   \ADIO27.PULLUP  (
    .O(ADIO27)
  );
  X_PU   \ADIO28.PULLUP  (
    .O(ADIO28)
  );
  X_PU   \ADIO29.PULLUP  (
    .O(ADIO29)
  );
  X_PU   \ADIO3.PULLUP  (
    .O(ADIO3)
  );
  X_PU   \ADIO30.PULLUP  (
    .O(ADIO30)
  );
  X_PU   \ADIO31.PULLUP  (
    .O(ADIO31)
  );
  X_PU   \ADIO32.PULLUP  (
    .O(ADIO32)
  );
  X_PU   \ADIO33.PULLUP  (
    .O(ADIO33)
  );
  X_PU   \ADIO34.PULLUP  (
    .O(ADIO34)
  );
  X_PU   \ADIO35.PULLUP  (
    .O(ADIO35)
  );
  X_PU   \ADIO36.PULLUP  (
    .O(ADIO36)
  );
  X_PU   \ADIO37.PULLUP  (
    .O(ADIO37)
  );
  X_PU   \ADIO38.PULLUP  (
    .O(ADIO38)
  );
  X_PU   \ADIO39.PULLUP  (
    .O(ADIO39)
  );
  X_PU   \ADIO4.PULLUP  (
    .O(ADIO4)
  );
  X_PU   \ADIO40.PULLUP  (
    .O(ADIO40)
  );
  X_PU   \ADIO41.PULLUP  (
    .O(ADIO41)
  );
  X_PU   \ADIO42.PULLUP  (
    .O(ADIO42)
  );
  X_PU   \ADIO43.PULLUP  (
    .O(ADIO43)
  );
  X_PU   \ADIO44.PULLUP  (
    .O(ADIO44)
  );
  X_PU   \ADIO45.PULLUP  (
    .O(ADIO45)
  );
  X_PU   \ADIO46.PULLUP  (
    .O(ADIO46)
  );
  X_PU   \ADIO47.PULLUP  (
    .O(ADIO47)
  );
  X_PU   \ADIO48.PULLUP  (
    .O(ADIO48)
  );
  X_PU   \ADIO49.PULLUP  (
    .O(ADIO49)
  );
  X_PU   \ADIO5.PULLUP  (
    .O(ADIO5)
  );
  X_PU   \ADIO50.PULLUP  (
    .O(ADIO50)
  );
  X_PU   \ADIO51.PULLUP  (
    .O(ADIO51)
  );
  X_PU   \ADIO52.PULLUP  (
    .O(ADIO52)
  );
  X_PU   \ADIO53.PULLUP  (
    .O(ADIO53)
  );
  X_PU   \ADIO54.PULLUP  (
    .O(ADIO54)
  );
  X_PU   \ADIO55.PULLUP  (
    .O(ADIO55)
  );
  X_PU   \ADIO56.PULLUP  (
    .O(ADIO56)
  );
  X_PU   \ADIO57.PULLUP  (
    .O(ADIO57)
  );
  X_PU   \ADIO58.PULLUP  (
    .O(ADIO58)
  );
  X_PU   \ADIO59.PULLUP  (
    .O(ADIO59)
  );
  X_PU   \ADIO6.PULLUP  (
    .O(ADIO6)
  );
  X_PU   \ADIO60.PULLUP  (
    .O(ADIO60)
  );
  X_PU   \ADIO61.PULLUP  (
    .O(ADIO61)
  );
  X_PU   \ADIO62.PULLUP  (
    .O(ADIO62)
  );
  X_PU   \ADIO63.PULLUP  (
    .O(ADIO63)
  );
  X_PU   \ADIO7.PULLUP  (
    .O(ADIO7)
  );
  X_PU   \ADIO8.PULLUP  (
    .O(ADIO8)
  );
  X_PU   \ADIO9.PULLUP  (
    .O(ADIO9)
  );
  X_AND4   \MASTER/$4I3271  (
    .I0(\NlwInverterSignal_MASTER/$4I3271/I0 ),
    .I1(\NlwInverterSignal_MASTER/$4I3271/I1 ),
    .I2(\NlwInverterSignal_MASTER/$4I3271/I2 ),
    .I3(SLOT64),
    .O(\MASTER/NS_IREAD64 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \MASTER/REQO_OE  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(CLK),
    .I(\MASTER/$4N3252 ),
    .O(OE_REQ),
    .RST(GND)
  );
  X_BUF   \MASTER/$4I3208  (
    .I(\MASTER/REG_0CH8 ),
    .O(\MASTER/LAT_TIME0 )
  );
  X_BUF   \MASTER/$4I3207  (
    .I(\MASTER/REG_0CH9 ),
    .O(\MASTER/LAT_TIME1 )
  );
  X_BUF   \MASTER/$4I3206  (
    .I(\MASTER/REG_0CH10 ),
    .O(\MASTER/LAT_TIME2 )
  );
  X_BUF   \MASTER/$4I3205  (
    .I(\MASTER/REG_0CH11 ),
    .O(\MASTER/LAT_TIME3 )
  );
  X_BUF   \MASTER/$4I3204  (
    .I(\MASTER/REG_0CH12 ),
    .O(\MASTER/LAT_TIME4 )
  );
  X_BUF   \MASTER/$4I3203  (
    .I(\MASTER/REG_0CH13 ),
    .O(\MASTER/LAT_TIME5 )
  );
  X_BUF   \MASTER/$4I3202  (
    .I(\MASTER/REG_0CH14 ),
    .O(\MASTER/LAT_TIME6 )
  );
  X_BUF   \MASTER/$4I3201  (
    .I(\MASTER/REG_0CH15 ),
    .O(\MASTER/LAT_TIME7 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \MASTER/$4I3116  (
    .CE(VCC),
    .CLK(CLK),
    .I(\MASTER/NS_IREAD64 ),
    .O(\MASTER/IREAD64 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND4   \MASTER/$4I3102  (
    .I0(\NlwInverterSignal_MASTER/$4I3102/I0 ),
    .I1(\NlwInverterSignal_MASTER/$4I3102/I1 ),
    .I2(\MASTER/IREAD64 ),
    .I3(M_DATA_INT),
    .O(IPWIN64)
  );
  X_AND2   \MASTER/$4I3072  (
    .I0(\NlwInverterSignal_MASTER/$4I3072/I0 ),
    .I1(\MASTER/DEV_TO ),
    .O(SET13)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \MASTER/$4I3068  (
    .CE(ADDR_BE),
    .CLK(CLK),
    .I(\MASTER/$4N3021 ),
    .O(\MASTER/$4N3030 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND3   \MASTER/$4I3051  (
    .I0(\NlwInverterSignal_MASTER/$4I3051/I0 ),
    .I1(\DEVSEL- ),
    .I2(M_DATA_INT),
    .O(SET12)
  );
  X_OR2   \MASTER/$4I2899  (
    .I0(M_ENABLE),
    .I1(CFG_SELF),
    .O(\MASTER/M_ENABLE )
  );
  X_AND4   \MASTER/$4I2686  (
    .I0(\NlwInverterSignal_MASTER/$4I2686/I0 ),
    .I1(\NlwInverterSignal_MASTER/$4I2686/I1 ),
    .I2(\NlwInverterSignal_MASTER/$4I2686/I2 ),
    .I3(M_DATA_INT),
    .O(IPWIN)
  );
  X_AND2   \MASTER/I_IDLE/$1I2807  (
    .I0(\NlwInverterSignal_MASTER/I_IDLE/$1I2807/I0 ),
    .I1(DR_BUS_INT),
    .O(\MASTER/I_IDLE/EQ-C )
  );
  X_AND2   \MASTER/I_IDLE/$1I2773  (
    .I0(\MASTER/M_ENABLE ),
    .I1(\MASTER/REQUEST ),
    .O(\MASTER/I_IDLE/VALIDREQ )
  );
  X_OR2   \MASTER/I_IDLE/$1I2770  (
    .I0(\GNT- ),
    .I1(\MASTER/I_IDLE/VALIDREQ ),
    .O(\MASTER/I_IDLE/$1N2776 )
  );
  X_AND4   \MASTER/I_IDLE/$1I2715  (
    .I0(\NlwInverterSignal_MASTER/I_IDLE/$1I2715/I0 ),
    .I1(\NlwInverterSignal_MASTER/I_IDLE/$1I2715/I1 ),
    .I2(\IRDY- ),
    .I3(\FRAME- ),
    .O(\NlwInverterSignal_MASTER/I_IDLE/$1I2715/O )
  );
  X_AND2   \MASTER/I_IDLE/$1I2698  (
    .I0(\MASTER/I_IDLE/ADDR_GNT ),
    .I1(I_IDLE_INT),
    .O(\MASTER/I_IDLE/I_IDLE_ADDR_GNT )
  );
  X_OR2   \MASTER/I_IDLE/$1I2647  (
    .I0(\NlwInverterSignal_MASTER/I_IDLE/$1I2647/I0 ),
    .I1(\MASTER/I_IDLE/PRE_C2 ),
    .O(\MASTER/I_IDLE/M_DATA_C2 )
  );
  X_AND2   \MASTER/I_IDLE/$1I2599  (
    .I0(\MASTER/I_IDLE/EQ-C ),
    .I1(\MASTER/I_IDLE/$1N2776 ),
    .O(\MASTER/I_IDLE/EQ-B )
  );
  X_OR2   \MASTER/I_IDLE/$1I2596  (
    .I0(\MASTER/I_IDLE/EQ-B ),
    .I1(\MASTER/I_IDLE/EQ-A ),
    .O(\MASTER/I_IDLE/M_DATA_AND_DR_BUS )
  );
  X_AND2   \MASTER/I_IDLE/$1I2595  (
    .I0(\GNT- ),
    .I1(M_DATA_INT),
    .O(\MASTER/I_IDLE/M_DATA_C1 )
  );
  X_AND4   \MASTER/I_IDLE/$1I2594  (
    .I0(\NlwInverterSignal_MASTER/I_IDLE/$1I2594/I0 ),
    .I1(\STOP- ),
    .I2(\TRDY- ),
    .I3(\MASTER/IFRAME- ),
    .O(\MASTER/I_IDLE/PRE_C2 )
  );
  X_AND2   \MASTER/I_IDLE/$1I2593  (
    .I0(\NlwInverterSignal_MASTER/I_IDLE/$1I2593/I0 ),
    .I1(\MASTER/I_IDLE/M_DATA_C1 ),
    .O(\MASTER/I_IDLE/EQ-A )
  );
  X_OR2   \MASTER/I_IDLE/$1I2592  (
    .I0(\MASTER/I_IDLE/I_IDLE_ADDR_GNT ),
    .I1(\MASTER/I_IDLE/M_DATA_AND_DR_BUS ),
    .O(\MASTER/I_IDLE/NS_I_IDLE )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \MASTER/I_IDLE/I_IDLE_FF  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(CLK),
    .I(\MASTER/I_IDLE/NS_I_IDLE ),
    .O(I_IDLE_INT),
    .RST(GND)
  );
  X_AND3   \MASTER/ADDR/$1I2632  (
    .I0(\NlwInverterSignal_MASTER/ADDR/$1I2632/I0 ),
    .I1(IRDY_M),
    .I2(FRAME_I),
    .O(\MASTER/ADDR/$1N2628 )
  );
  X_AND2   \MASTER/ADDR/$1I2630  (
    .I0(\MASTER/ADDR/M_ADDR_DEAD ),
    .I1(\MASTER/ADDR/$1N2628 ),
    .O(\NlwInverterSignal_MASTER/ADDR/$1I2630/O )
  );
  X_AND3   \MASTER/ADDR/$1I2623  (
    .I0(\NlwInverterSignal_MASTER/ADDR/$1I2623/I0 ),
    .I1(\MASTER/M_ENABLE ),
    .I2(\MASTER/REQUEST ),
    .O(\MASTER/ADDR/M_ADDR_DEAD )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \MASTER/ADDR/MAN_FF  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(CLK),
    .I(\MASTER/ADDR/NS_MAN ),
    .O(M_ADDR_N),
    .RST(GND)
  );
  X_AND3   \MASTER/ADDR/$1I2602  (
    .I0(\NlwInverterSignal_MASTER/ADDR/$1I2602/I0 ),
    .I1(IRDY_M),
    .I2(FRAME_I),
    .O(\MASTER/ADDR/$1N2603 )
  );
  X_AND2   \MASTER/ADDR/$1I2599  (
    .I0(\MASTER/ADDR/M_ADDR_DEAD ),
    .I1(\MASTER/ADDR/$1N2603 ),
    .O(\MASTER/ADDR/NS_ABE )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \MASTER/ADDR/ABE_FF  (
    .CE(VCC),
    .CLK(CLK),
    .I(\MASTER/ADDR/NS_ABE ),
    .O(ADDR_BE),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND4   \MASTER/DR_BUS/$1I2913  (
    .I0(\NlwInverterSignal_MASTER/DR_BUS/$1I2913/I0 ),
    .I1(\NlwInverterSignal_MASTER/DR_BUS/$1I2913/I1 ),
    .I2(\NlwInverterSignal_MASTER/DR_BUS/$1I2913/I2 ),
    .I3(I_IDLE_INT),
    .O(\MASTER/DR_BUS/EQN-B0 )
  );
  X_OR2   \MASTER/DR_BUS/$1I2819  (
    .I0(\MASTER/DR_BUS/$1N2820 ),
    .I1(\MASTER/DR_BUS/COMMON-A ),
    .O(\MASTER/DR_BUS/EQN-A1 )
  );
  X_AND2   \MASTER/DR_BUS/$1I2808  (
    .I0(\MASTER/DR_BUS/$1N2812 ),
    .I1(DR_BUS_INT),
    .O(\MASTER/DR_BUS/COMMON-B )
  );
  X_OR2   \MASTER/DR_BUS/$1I2805  (
    .I0(\NlwInverterSignal_MASTER/DR_BUS/$1I2805/I0 ),
    .I1(\NlwInverterSignal_MASTER/DR_BUS/$1I2805/I1 ),
    .O(\MASTER/DR_BUS/$1N2812 )
  );
  X_OR2   \MASTER/DR_BUS/$1I2789  (
    .I0(\MASTER/DR_BUS/$1N2793 ),
    .I1(\MASTER/DR_BUS/COMMON-A ),
    .O(\MASTER/DR_BUS/EQN-A0 )
  );
  X_AND2   \MASTER/DR_BUS/$1I2787  (
    .I0(\NlwInverterSignal_MASTER/DR_BUS/$1I2787/I0 ),
    .I1(\MASTER/DR_BUS/AAARGH ),
    .O(\MASTER/DR_BUS/$1N2820 )
  );
  X_AND3   \MASTER/DR_BUS/$1I2757  (
    .I0(\IRDY- ),
    .I1(\FRAME- ),
    .I2(\MASTER/DR_BUS/EQN-B1 ),
    .O(\MASTER/DR_BUS/$1N2745 )
  );
  X_AND3   \MASTER/DR_BUS/$1I2752  (
    .I0(\NlwInverterSignal_MASTER/DR_BUS/$1I2752/I0 ),
    .I1(\NlwInverterSignal_MASTER/DR_BUS/$1I2752/I1 ),
    .I2(I_IDLE_INT),
    .O(\MASTER/DR_BUS/EQN-B1 )
  );
  X_OR2   \MASTER/DR_BUS/$1I2744  (
    .I0(\MASTER/DR_BUS/$1N2745 ),
    .I1(\MASTER/DR_BUS/EQN-A1 ),
    .O(\MASTER/DR_BUS/NS_1 )
  );
  X_AND3   \MASTER/DR_BUS/$1I2732  (
    .I0(\NlwInverterSignal_MASTER/DR_BUS/$1I2732/I0 ),
    .I1(\NlwInverterSignal_MASTER/DR_BUS/$1I2732/I1 ),
    .I2(\MASTER/DR_BUS/COMMON-B ),
    .O(\MASTER/DR_BUS/$1N2793 )
  );
  X_AND2   \MASTER/DR_BUS/$1I2721  (
    .I0(\NlwInverterSignal_MASTER/DR_BUS/$1I2721/I0 ),
    .I1(\MASTER/DR_BUS/$1N2720 ),
    .O(\MASTER/DR_BUS/COMMON-A )
  );
  X_OR2   \MASTER/DR_BUS/$1I2719  (
    .I0(\NlwInverterSignal_MASTER/DR_BUS/$1I2719/I0 ),
    .I1(\MASTER/DR_BUS/$1N2718 ),
    .O(\MASTER/DR_BUS/COND )
  );
  X_AND3   \MASTER/DR_BUS/$1I2712  (
    .I0(\FRAME- ),
    .I1(\IRDY- ),
    .I2(\MASTER/DR_BUS/EQN-B0 ),
    .O(\MASTER/DR_BUS/$1N2700 )
  );
  X_AND4   \MASTER/DR_BUS/$1I2706  (
    .I0(\NlwInverterSignal_MASTER/DR_BUS/$1I2706/I0 ),
    .I1(\STOP- ),
    .I2(\TRDY- ),
    .I3(\MASTER/IFRAME- ),
    .O(\MASTER/DR_BUS/$1N2718 )
  );
  X_AND2   \MASTER/DR_BUS/$1I2704  (
    .I0(\NlwInverterSignal_MASTER/DR_BUS/$1I2704/I0 ),
    .I1(M_DATA_INT),
    .O(\MASTER/DR_BUS/$1N2720 )
  );
  X_OR2   \MASTER/DR_BUS/$1I2699  (
    .I0(\MASTER/DR_BUS/$1N2700 ),
    .I1(\MASTER/DR_BUS/EQN-A0 ),
    .O(\MASTER/DR_BUS/NS_0 )
  );
  X_MUX2   \MASTER/DR_BUS/$1I2498  (
    .IA(\MASTER/DR_BUS/NS_0 ),
    .IB(\MASTER/DR_BUS/NS_1 ),
    .O(\MASTER/DR_BUS/NS_DR_BUS ),
    .SEL(GNT_IN)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \MASTER/DR_BUS/DR_BUS_FF  (
    .CE(VCC),
    .CLK(CLK),
    .I(\MASTER/DR_BUS/NS_DR_BUS ),
    .O(DR_BUS_INT),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND2   \MASTER/DR_BUS/$1I2908/$1I9  (
    .I0(DR_BUS_INT),
    .I1(\$1N4834 ),
    .O(\MASTER/DR_BUS/$1I2908/M1 )
  );
  X_OR2   \MASTER/DR_BUS/$1I2908/$1I8  (
    .I0(\MASTER/DR_BUS/$1I2908/M1 ),
    .I1(\MASTER/DR_BUS/$1I2908/M0 ),
    .O(\MASTER/DR_BUS/AAARGH )
  );
  X_AND2   \MASTER/DR_BUS/$1I2908/$1I7  (
    .I0(\NlwInverterSignal_MASTER/DR_BUS/$1I2908/$1I7/I0 ),
    .I1(\MASTER/DR_BUS/COMMON-B ),
    .O(\MASTER/DR_BUS/$1I2908/M0 )
  );
  X_AND2   \MASTER/DR_BUS/$1I2917/$1I9  (
    .I0(\MASTER/DR_BUS/$1N2925 ),
    .I1(\$1N4834 ),
    .O(\MASTER/DR_BUS/$1I2917/M1 )
  );
  X_OR2   \MASTER/DR_BUS/$1I2917/$1I8  (
    .I0(\MASTER/DR_BUS/$1I2917/M1 ),
    .I1(\MASTER/DR_BUS/$1I2917/M0 ),
    .O(\MASTER/DR_BUS/BBBRGH )
  );
  X_AND2   \MASTER/DR_BUS/$1I2917/$1I7  (
    .I0(\NlwInverterSignal_MASTER/DR_BUS/$1I2917/$1I7/I0 ),
    .I1(\MASTER/REQUEST ),
    .O(\MASTER/DR_BUS/$1I2917/M0 )
  );
  X_ZERO   \MASTER/DR_BUS/$1I2927/$1I2218  (
    .O(\MASTER/DR_BUS/$1I2927/$1N2216 )
  );
  X_BUF   \MASTER/DR_BUS/$1I2927/L  (
    .I(\MASTER/DR_BUS/$1I2927/$1N2216 ),
    .O(\MASTER/DR_BUS/$1N2925 )
  );
  X_AND2   \MASTER/M_DATA/$1I2590  (
    .I0(\NlwInverterSignal_MASTER/M_DATA/$1I2590/I0 ),
    .I1(ADDR_BE),
    .O(\MASTER/M_DATA/EQN_B )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \MASTER/M_DATA/M_DATA1  (
    .CE(VCC),
    .CLK(CLK),
    .I(\MASTER/M_DATA/NS_MDATA ),
    .O(M_DATA),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_OR2   \MASTER/M_DATA/$1I2518  (
    .I0(\NlwInverterSignal_MASTER/M_DATA/$1I2518/I0 ),
    .I1(\MASTER/M_DATA/$1N2519 ),
    .O(\MASTER/M_DATA/EQN-A )
  );
  X_AND4   \MASTER/M_DATA/$1I2502  (
    .I0(\NlwInverterSignal_MASTER/M_DATA/$1I2502/I0 ),
    .I1(\STOP- ),
    .I2(\TRDY- ),
    .I3(\MASTER/IFRAME- ),
    .O(\MASTER/M_DATA/$1N2519 )
  );
  X_AND2   \MASTER/M_DATA/$1I2499  (
    .I0(\MASTER/M_DATA/EQN-A ),
    .I1(M_DATA_INT),
    .O(\MASTER/M_DATA/$1N2507 )
  );
  X_OR2   \MASTER/M_DATA/$1I2498  (
    .I0(\MASTER/M_DATA/$1N2507 ),
    .I1(\MASTER/M_DATA/EQN_B ),
    .O(\MASTER/M_DATA/NS_MDATA )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \MASTER/M_DATA/M_DATA  (
    .CE(VCC),
    .CLK(CLK),
    .I(\MASTER/M_DATA/NS_MDATA ),
    .O(M_DATA_INT),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_OR2   \MASTER/$1I2914/$1I2956  (
    .I0(MIKELOVEJOY),
    .I1(\MASTER/$1I2914/$1N2959 ),
    .O(\MASTER/$1I2914/END_OF_XFER )
  );
  X_OR2   \MASTER/$1I2914/$1I2952  (
    .I0(MIKELOVEJOY),
    .I1(ADDR_BE),
    .O(\MASTER/$1I2914/CANCEL )
  );
  X_OR3   \MASTER/$1I2914/$1I2947  (
    .I0(\NlwInverterSignal_MASTER/$1I2914/$1I2947/I0 ),
    .I1(\MASTER/REQUEST ),
    .I2(EX),
    .O(\MASTER/$1I2914/LOCKOUT )
  );
  X_AND2   \MASTER/$1I2914/$1I2931  (
    .I0(\NlwInverterSignal_MASTER/$1I2914/$1I2931/I0 ),
    .I1(\MASTER/$1I2914/$1N2938 ),
    .O(\MASTER/$1I2914/$1N2929 )
  );
  X_OR2   \MASTER/$1I2914/$1I2930  (
    .I0(\MASTER/$1I2914/SCG64 ),
    .I1(REQUEST64),
    .O(\MASTER/$1I2914/$1N2938 )
  );
  X_AND2   \MASTER/$1I2914/$1I2927  (
    .I0(\NlwInverterSignal_MASTER/$1I2914/$1I2927/I0 ),
    .I1(\MASTER/$1I2914/M_DATA_Q ),
    .O(\MASTER/$1I2914/$1N2959 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \MASTER/$1I2914/$1I2926  (
    .CE(VCC),
    .CLK(CLK),
    .I(M_DATA_INT),
    .O(\MASTER/$1I2914/M_DATA_Q ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND3   \MASTER/$1I2914/$1I2908  (
    .I0(\NlwInverterSignal_MASTER/$1I2914/$1I2908/I0 ),
    .I1(\MASTER/$1I2914/ADDR_BE_Q ),
    .I2(\MASTER/$1I2914/REQUEST64Q ),
    .O(\MASTER/$1I2914/SCG64 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \MASTER/$1I2914/$1I2903  (
    .CE(VCC),
    .CLK(CLK),
    .I(\MASTER/REQUEST64 ),
    .O(\MASTER/$1I2914/REQUEST64Q ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND2   \MASTER/$1I2914/$1I2895  (
    .I0(\NlwInverterSignal_MASTER/$1I2914/$1I2895/I0 ),
    .I1(\MASTER/$1I2914/$1N2897 ),
    .O(\MASTER/$1I2914/$1N2894 )
  );
  X_OR2   \MASTER/$1I2914/$1I2893  (
    .I0(\MASTER/$1I2914/SCG64 ),
    .I1(REQUEST64),
    .O(\MASTER/$1I2914/$1N2897 )
  );
  X_AND2   \MASTER/$1I2914/$1I2880  (
    .I0(\NlwInverterSignal_MASTER/$1I2914/$1I2880/I0 ),
    .I1(\MASTER/$1I2914/ADDR_BE_Q ),
    .O(\MASTER/$1I2914/SCG32 )
  );
  X_AND2   \MASTER/$1I2914/$1I2879  (
    .I0(\NlwInverterSignal_MASTER/$1I2914/$1I2879/I0 ),
    .I1(\MASTER/$1I2914/$1N2884 ),
    .O(\MASTER/$1I2914/$1N2881 )
  );
  X_OR4   \MASTER/$1I2914/$1I2878  (
    .I0(\MASTER/$1I2914/SCG64 ),
    .I1(\MASTER/$1I2914/SCG32 ),
    .I2(REQUEST64),
    .I3(REQUEST),
    .O(\MASTER/$1I2914/$1N2884 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \MASTER/$1I2914/$1I2862  (
    .CE(VCC),
    .CLK(CLK),
    .I(ADDR_BE),
    .O(\MASTER/$1I2914/ADDR_BE_Q ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_OR2   \MASTER/$1I2914/$1I2853/$1I2214  (
    .I0(\MASTER/$1I2914/$1N2881 ),
    .I1(\MASTER/REQUEST ),
    .O(\MASTER/$1I2914/$1I2853/$1N2215 )
  );
  X_AND2   \MASTER/$1I2914/$1I2853/$1I2213  (
    .I0(\NlwInverterSignal_MASTER/$1I2914/$1I2853/$1I2213/I0 ),
    .I1(\MASTER/$1I2914/$1I2853/$1N2215 ),
    .O(\MASTER/$1I2914/$1I2853/D )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \MASTER/$1I2914/$1I2853/FDCE  (
    .CE(VCC),
    .CLK(CLK),
    .I(\MASTER/$1I2914/$1I2853/D ),
    .O(\MASTER/REQUEST ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_OR2   \MASTER/$1I2914/$1I2864/$1I2214  (
    .I0(\MASTER/$1I2914/$1N2894 ),
    .I1(\MASTER/REQUEST64 ),
    .O(\MASTER/$1I2914/$1I2864/$1N2215 )
  );
  X_AND2   \MASTER/$1I2914/$1I2864/$1I2213  (
    .I0(\NlwInverterSignal_MASTER/$1I2914/$1I2864/$1I2213/I0 ),
    .I1(\MASTER/$1I2914/$1I2864/$1N2215 ),
    .O(\MASTER/$1I2914/$1I2864/D )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \MASTER/$1I2914/$1I2864/FDCE  (
    .CE(VCC),
    .CLK(CLK),
    .I(\MASTER/$1I2914/$1I2864/D ),
    .O(\MASTER/REQUEST64 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_OR2   \MASTER/$1I2914/$1I2932/$1I2214  (
    .I0(\MASTER/$1I2914/$1N2929 ),
    .I1(ATTEMPT64),
    .O(\MASTER/$1I2914/$1I2932/$1N2215 )
  );
  X_AND2   \MASTER/$1I2914/$1I2932/$1I2213  (
    .I0(\NlwInverterSignal_MASTER/$1I2914/$1I2932/$1I2213/I0 ),
    .I1(\MASTER/$1I2914/$1I2932/$1N2215 ),
    .O(\MASTER/$1I2914/$1I2932/D )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \MASTER/$1I2914/$1I2932/FDCE  (
    .CE(VCC),
    .CLK(CLK),
    .I(\MASTER/$1I2914/$1I2932/D ),
    .O(ATTEMPT64),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND2   \MASTER/FRAME/$2I3529  (
    .I0(\MASTER/FRAME/DTO ),
    .I1(NlwRenamedSig_OI_TIME_OUT),
    .O(\MASTER/FRAME/$2N3531 )
  );
  X_OR3   \MASTER/FRAME/$2I3528  (
    .I0(\NlwInverterSignal_MASTER/FRAME/$2I3528/I0 ),
    .I1(COMPLETE),
    .I2(\MASTER/FRAME/$2N3531 ),
    .O(\MASTER/FRAME/DONE_1 )
  );
  X_AND2   \MASTER/FRAME/$2I3518  (
    .I0(\MASTER/FRAME/DTO ),
    .I1(NlwRenamedSig_OI_TIME_OUT),
    .O(\MASTER/FRAME/$2N3521 )
  );
  X_OR3   \MASTER/FRAME/$2I3511  (
    .I0(\NlwInverterSignal_MASTER/FRAME/$2I3511/I0 ),
    .I1(COMPLETE),
    .I2(\MASTER/FRAME/$2N3521 ),
    .O(\MASTER/FRAME/DONE_0 )
  );
  X_OR2   \MASTER/FRAME/$2I3495  (
    .I0(\IIRDY_I- ),
    .I1(\MASTER/IFRAME- ),
    .O(\MASTER/FRAME/INITIAL )
  );
  X_AND2   \MASTER/FRAME/$2I3468  (
    .I0(M_READY),
    .I1(\MASTER/FRAME/DONE_0 ),
    .O(\MASTER/FRAME/$2N3475 )
  );
  X_AND2   \MASTER/FRAME/$2I3464  (
    .I0(\NlwInverterSignal_MASTER/FRAME/$2I3464/I0 ),
    .I1(\MASTER/FRAME/FEEDBACK ),
    .O(\MASTER/FRAME/KO_T_0 )
  );
  X_AND2   \MASTER/FRAME/$2I3463  (
    .I0(\NlwInverterSignal_MASTER/FRAME/$2I3463/I0 ),
    .I1(\MASTER/FRAME/FEEDBACK ),
    .O(\MASTER/FRAME/KO_T_1 )
  );
  X_AND2   \MASTER/FRAME/$2I3459  (
    .I0(M_READY),
    .I1(\MASTER/FRAME/$2N3450 ),
    .O(\MASTER/FRAME/$2N3449 )
  );
  X_AND2   \MASTER/FRAME/$2I3458  (
    .I0(\MASTER/FRAME/INITIAL ),
    .I1(\MASTER/FRAME/DONE_1 ),
    .O(\MASTER/FRAME/$2N3450 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \MASTER/FRAME/IFRAME_I-  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(FRAME_CE),
    .CLK(CLK),
    .I(\NS_FRAME- ),
    .O(\IFRAME_I- ),
    .RST(GND)
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \MASTER/FRAME/IFRAME-  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(CLK),
    .I(\IFRAME_I- ),
    .O(\MASTER/IFRAME- ),
    .RST(GND)
  );
  X_OR2   \MASTER/FRAME/$1I3470  (
    .I0(\MASTER/FRAME/TURN_ON ),
    .I1(\MASTER/FRAME/$1N3468 ),
    .O(\NlwInverterSignal_MASTER/FRAME/$1I3470/O )
  );
  X_AND2   \MASTER/FRAME/$1I3466  (
    .I0(\NlwInverterSignal_MASTER/FRAME/$1I3466/I0 ),
    .I1(ADDR_BE),
    .O(\MASTER/FRAME/TURN_ON )
  );
  X_MUX2   \MASTER/FRAME/$1I3419  (
    .IA(\MASTER/FRAME/NS_S_0 ),
    .IB(\MASTER/FRAME/NS_S_1 ),
    .O(\NS_FRAME- ),
    .SEL(STOP_I)
  );
  X_AND2   \MASTER/FRAME/$1I3393  (
    .I0(\NlwInverterSignal_MASTER/FRAME/$1I3393/I0 ),
    .I1(\MASTER/FRAME/FEEDBACK ),
    .O(\MASTER/FRAME/$1N3369 )
  );
  X_OR2   \MASTER/FRAME/$1I3368  (
    .I0(\MASTER/FRAME/TURN_ON ),
    .I1(\MASTER/FRAME/$1N3369 ),
    .O(\NlwInverterSignal_MASTER/FRAME/$1I3368/O )
  );
  X_AND4   \MASTER/FRAME/$1I3323  (
    .I0(\NlwInverterSignal_MASTER/FRAME/$1I3323/I0 ),
    .I1(STOP_I),
    .I2(ACK64_I),
    .I3(\MASTER/FRAME/IRDY_64 ),
    .O(\NlwInverterSignal_MASTER/FRAME/$1I3323/O )
  );
  X_AND2   \MASTER/FRAME/$1I3322  (
    .I0(\NlwInverterSignal_MASTER/FRAME/$1I3322/I0 ),
    .I1(ATTEMPT64),
    .O(\MASTER/FRAME/IRDY_64 )
  );
  X_AND4   \MASTER/FRAME/$1I3144  (
    .I0(\NlwInverterSignal_MASTER/FRAME/$1I3144/I0 ),
    .I1(\NlwInverterSignal_MASTER/FRAME/$1I3144/I1 ),
    .I2(\NlwInverterSignal_MASTER/FRAME/$1I3144/I2 ),
    .I3(M_DATA_INT),
    .O(\MASTER/FRAME/FEEDBACK )
  );
  X_BUF   \MASTER/FRAME/$1I2554/NC  (
    .I(\MASTER/REQUEST ),
    .O(\NLW_MASTER/FRAME/$1I2554/NC_O_UNCONNECTED )
  );
  X_AND2   \MASTER/FRAME/$1I3467/$1I9  (
    .I0(\MASTER/FRAME/KO_T_1 ),
    .I1(TRDY_M),
    .O(\MASTER/FRAME/$1I3467/M1 )
  );
  X_OR2   \MASTER/FRAME/$1I3467/$1I8  (
    .I0(\MASTER/FRAME/$1I3467/M1 ),
    .I1(\MASTER/FRAME/$1I3467/M0 ),
    .O(\MASTER/FRAME/$1N3468 )
  );
  X_AND2   \MASTER/FRAME/$1I3467/$1I7  (
    .I0(\NlwInverterSignal_MASTER/FRAME/$1I3467/$1I7/I0 ),
    .I1(\MASTER/FRAME/KO_T_0 ),
    .O(\MASTER/FRAME/$1I3467/M0 )
  );
  X_AND2   \MASTER/FRAME/$2I3559/$1I9  (
    .I0(GNT_IN),
    .I1(CFG254),
    .O(\MASTER/FRAME/$2I3559/M1 )
  );
  X_OR2   \MASTER/FRAME/$2I3559/$1I8  (
    .I0(\MASTER/FRAME/$2I3559/M1 ),
    .I1(\MASTER/FRAME/$2I3559/M0 ),
    .O(\MASTER/FRAME/DTO )
  );
  X_AND2   \MASTER/FRAME/$2I3559/$1I7  (
    .I0(\NlwInverterSignal_MASTER/FRAME/$2I3559/$1I7/I0 ),
    .I1(\GNT- ),
    .O(\MASTER/FRAME/$2I3559/M0 )
  );
  X_AND2   \MASTER/IRDY/$2I3437  (
    .I0(\NlwInverterSignal_MASTER/IRDY/$2I3437/I0 ),
    .I1(M_DATA_INT),
    .O(\MASTER/IRDY/EQN-F )
  );
  X_AND3   \MASTER/IRDY/$2I3435  (
    .I0(\MASTER/IRDY/EQN-E ),
    .I1(M_READY),
    .I2(\MASTER/IRDY/EQN-F ),
    .O(\NlwInverterSignal_MASTER/IRDY/$2I3435/O )
  );
  X_AND2   \MASTER/IRDY/$2I3390  (
    .I0(\MASTER/IRDY/$2N3294 ),
    .I1(\MASTER/IRDY/ALLOWED ),
    .O(\NlwInverterSignal_MASTER/IRDY/$2I3390/O )
  );
  X_AND2   \MASTER/IRDY/$2I3387  (
    .I0(\MASTER/IRDY/$2N3385 ),
    .I1(M_FIRST),
    .O(\MASTER/IRDY/M_FIRST1 )
  );
  X_OR2   \MASTER/IRDY/$2I3380  (
    .I0(\MASTER/IRDY/END_OF_INIT ),
    .I1(\MASTER/IRDY/$2N3383 ),
    .O(\MASTER/IRDY/M_FIRSTIN )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \MASTER/IRDY/M1FF  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(CLK),
    .I(\MASTER/IRDY/M_FIRSTIN ),
    .O(M_FIRST),
    .RST(GND)
  );
  X_AND2   \MASTER/IRDY/$2I3334  (
    .I0(M_FIRST),
    .I1(\MASTER/IRDY/$2N3355 ),
    .O(\MASTER/IRDY/M_FIRST0 )
  );
  X_AND2   \MASTER/IRDY/$2I3332  (
    .I0(\NlwInverterSignal_MASTER/IRDY/$2I3332/I0 ),
    .I1(\MASTER/IRDY/WS_A_0 ),
    .O(\NlwInverterSignal_MASTER/IRDY/$2I3332/O )
  );
  X_AND2   \MASTER/IRDY/$2I3233  (
    .I0(\NlwInverterSignal_MASTER/IRDY/$2I3233/I0 ),
    .I1(\MASTER/IRDY/M_DATA_Q ),
    .O(\MASTER/IRDY/END_OF_INIT )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \MASTER/IRDY/$2I3082  (
    .CE(VCC),
    .CLK(CLK),
    .I(M_DATA_INT),
    .O(\MASTER/IRDY/M_DATA_Q ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND4   \MASTER/IRDY/$1I3779  (
    .I0(\NlwInverterSignal_MASTER/IRDY/$1I3779/I0 ),
    .I1(M_READY),
    .I2(M_DATA_INT),
    .I3(\MASTER/IRDY/EQN-E ),
    .O(\NlwInverterSignal_MASTER/IRDY/$1I3779/O )
  );
  X_AND2   \MASTER/IRDY/$1I3742  (
    .I0(\MASTER/IRDY/EQN-E ),
    .I1(M_DATA_INT),
    .O(\MASTER/IRDY/$1N3756 )
  );
  X_OR2   \MASTER/IRDY/$1I3738  (
    .I0(\NlwInverterSignal_MASTER/IRDY/$1I3738/I0 ),
    .I1(\NlwInverterSignal_MASTER/IRDY/$1I3738/I1 ),
    .O(\MASTER/IRDY/EQN-G )
  );
  X_AND2   \MASTER/IRDY/$1I3735  (
    .I0(\MASTER/IRDY/EQN-G ),
    .I1(\MASTER/IRDY/$1N3756 ),
    .O(\MASTER/IRDY/$1N3772 )
  );
  X_AND2   \MASTER/IRDY/$1I3734  (
    .I0(\MASTER/IRDY/$1N3772 ),
    .I1(M_READY),
    .O(\MASTER/IRDY/ALLOWED )
  );
  X_OR2   \MASTER/IRDY/$1I3699  (
    .I0(\NlwInverterSignal_MASTER/IRDY/$1I3699/I0 ),
    .I1(\MASTER/IRDY/$1N3721 ),
    .O(\MASTER/IRDY/EQN-E )
  );
  X_AND3   \MASTER/IRDY/$1I3698  (
    .I0(\NlwInverterSignal_MASTER/IRDY/$1I3698/I0 ),
    .I1(\STOP- ),
    .I2(\TRDY- ),
    .O(\MASTER/IRDY/$1N3721 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \MASTER/IRDY/IIRDY-  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(CLK),
    .I(\IIRDY_I- ),
    .O(\MASTER/IIRDY- ),
    .RST(GND)
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \MASTER/IRDY/IIRDY_I-  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(IRDY_CE),
    .CLK(CLK),
    .I(\NS_IRDY- ),
    .O(\IIRDY_I- ),
    .RST(GND)
  );
  X_AND2   \MASTER/IRDY/$1I3498  (
    .I0(\NlwInverterSignal_MASTER/IRDY/$1I3498/I0 ),
    .I1(\MASTER/IRDY/$1N3502 ),
    .O(\MASTER/IRDY/WS_A_1 )
  );
  X_OR2   \MASTER/IRDY/$1I3497  (
    .I0(\IFRAME_I- ),
    .I1(ATTEMPT64),
    .O(\MASTER/IRDY/$1N3502 )
  );
  X_AND2   \MASTER/IRDY/$1I3491  (
    .I0(\NlwInverterSignal_MASTER/IRDY/$1I3491/I0 ),
    .I1(\IFRAME_I- ),
    .O(\MASTER/IRDY/WS_A_0 )
  );
  X_AND2   \MASTER/IRDY/$1I3487  (
    .I0(\NlwInverterSignal_MASTER/IRDY/$1I3487/I0 ),
    .I1(\MASTER/IRDY/$1N3493 ),
    .O(\NlwInverterSignal_MASTER/IRDY/$1I3487/O )
  );
  X_AND2   \MASTER/IRDY/$1I3211  (
    .I0(\MASTER/IRDY/CORE_READY ),
    .I1(\MASTER/IRDY/ALLOWED ),
    .O(\NlwInverterSignal_MASTER/IRDY/$1I3211/O )
  );
  X_AND2   \MASTER/IRDY/$1I3227/$1I9  (
    .I0(\MASTER/IRDY/NS_1 ),
    .I1(STOP_I),
    .O(\MASTER/IRDY/$1I3227/M1 )
  );
  X_OR2   \MASTER/IRDY/$1I3227/$1I8  (
    .I0(\MASTER/IRDY/$1I3227/M1 ),
    .I1(\MASTER/IRDY/$1I3227/M0 ),
    .O(\NS_IRDY- )
  );
  X_AND2   \MASTER/IRDY/$1I3227/$1I7  (
    .I0(\NlwInverterSignal_MASTER/IRDY/$1I3227/$1I7/I0 ),
    .I1(\MASTER/IRDY/NS_0 ),
    .O(\MASTER/IRDY/$1I3227/M0 )
  );
  X_AND2   \MASTER/IRDY/$1I3492/$1I9  (
    .I0(\MASTER/IRDY/WS_A_1 ),
    .I1(ACK64_I),
    .O(\MASTER/IRDY/$1I3492/M1 )
  );
  X_OR2   \MASTER/IRDY/$1I3492/$1I8  (
    .I0(\MASTER/IRDY/$1I3492/M1 ),
    .I1(\MASTER/IRDY/$1I3492/M0 ),
    .O(\MASTER/IRDY/$1N3493 )
  );
  X_AND2   \MASTER/IRDY/$1I3492/$1I7  (
    .I0(\NlwInverterSignal_MASTER/IRDY/$1I3492/$1I7/I0 ),
    .I1(\MASTER/IRDY/WS_A_0 ),
    .O(\MASTER/IRDY/$1I3492/M0 )
  );
  X_ONE   \MASTER/IRDY/$1I3563/$1I2220  (
    .O(\MASTER/IRDY/$1I3563/$1N2216 )
  );
  X_BUF   \MASTER/IRDY/$1I3563/H  (
    .I(\MASTER/IRDY/$1I3563/$1N2216 ),
    .O(IRDY_CE)
  );
  X_AND2   \MASTER/IRDY/$2I3285/$1I9  (
    .I0(\MASTER/IRDY/M_FIRST1 ),
    .I1(STOP_I),
    .O(\MASTER/IRDY/$2I3285/M1 )
  );
  X_OR2   \MASTER/IRDY/$2I3285/$1I8  (
    .I0(\MASTER/IRDY/$2I3285/M1 ),
    .I1(\MASTER/IRDY/$2I3285/M0 ),
    .O(\MASTER/IRDY/$2N3383 )
  );
  X_AND2   \MASTER/IRDY/$2I3285/$1I7  (
    .I0(\NlwInverterSignal_MASTER/IRDY/$2I3285/$1I7/I0 ),
    .I1(\MASTER/IRDY/M_FIRST0 ),
    .O(\MASTER/IRDY/$2I3285/M0 )
  );
  X_OR2   \MASTER/REQ/$1I2735  (
    .I0(MIKELOVEJOY),
    .I1(\MASTER/REQ/$1N2737 ),
    .O(\MASTER/REQ/SOXFER )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \MASTER/REQ/$1I2734  (
    .CE(VCC),
    .CLK(CLK),
    .I(\MASTER/S_TAR ),
    .O(\MASTER/REQ/S_TARQ ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_OR2   \MASTER/REQ/$1I2729  (
    .I0(\MASTER/REQ/NORM1 ),
    .I1(\MASTER/REQ/EXT ),
    .O(\MASTER/REQ/Y )
  );
  X_AND2   \MASTER/REQ/$1I2728  (
    .I0(\MASTER/REQUEST ),
    .I1(\MASTER/M_ENABLE ),
    .O(\MASTER/REQ/NORM2 )
  );
  X_OR2   \MASTER/REQ/$1I2726  (
    .I0(\MASTER/REQ/S_TARQ ),
    .I1(\MASTER/S_TAR ),
    .O(\NlwInverterSignal_MASTER/REQ/$1I2726/O )
  );
  X_AND2   \MASTER/REQ/$1I2722  (
    .I0(\MASTER/M_ENABLE ),
    .I1(REQUESTHOLD),
    .O(\MASTER/REQ/EXT )
  );
  X_AND2   \MASTER/REQ/$1I2721  (
    .I0(\MASTER/REQ/S_TAR_OR ),
    .I1(\MASTER/REQ/REQ_BUS ),
    .O(\NlwInverterSignal_MASTER/REQ/$1I2721/O )
  );
  X_AND2   \MASTER/REQ/$1I2719  (
    .I0(\MASTER/M_ENABLE ),
    .I1(\MASTER/REQUEST ),
    .O(\MASTER/REQ/NORM1 )
  );
  X_OR2   \MASTER/REQ/$1I2707  (
    .I0(\MASTER/REQ/X ),
    .I1(\MASTER/REQ/Y ),
    .O(\MASTER/REQ/REQ_BUS )
  );
  X_AND2   \MASTER/REQ/$1I2670  (
    .I0(\NlwInverterSignal_MASTER/REQ/$1I2670/I0 ),
    .I1(M_DATA_INT),
    .O(\MASTER/REQ/$1N2737 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \MASTER/REQ/$1I2669  (
    .CLK(CLK),
    .I(M_DATA_INT),
    .O(\MASTER/REQ/M_DATA_Q ),
    .RST(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \MASTER/REQ/IREQ-  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(CLK),
    .I(\MASTER/IREQ_I- ),
    .O(\MASTER/IREQ- ),
    .RST(GND)
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \MASTER/REQ/IREQ_I-  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(CLK),
    .I(\MASTER/NS_REQ- ),
    .O(\MASTER/IREQ_I- ),
    .RST(GND)
  );
  X_OR2   \MASTER/REQ/$1I2708/$1I2214  (
    .I0(\MASTER/REQ/NORM2 ),
    .I1(\MASTER/REQ/X ),
    .O(\MASTER/REQ/$1I2708/$1N2215 )
  );
  X_AND2   \MASTER/REQ/$1I2708/$1I2213  (
    .I0(\NlwInverterSignal_MASTER/REQ/$1I2708/$1I2213/I0 ),
    .I1(\MASTER/REQ/$1I2708/$1N2215 ),
    .O(\MASTER/REQ/$1I2708/D )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \MASTER/REQ/$1I2708/FDCE  (
    .CE(VCC),
    .CLK(CLK),
    .I(\MASTER/REQ/$1I2708/D ),
    .O(\MASTER/REQ/X ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND2   \MASTER/REQ64/$2I3435  (
    .I0(M_READY),
    .I1(\MASTER/REQ64/DONE_0 ),
    .O(\MASTER/REQ64/$2N3428 )
  );
  X_AND2   \MASTER/REQ64/$2I3432  (
    .I0(\MASTER/REQ64/INITIAL ),
    .I1(\MASTER/REQ64/DONE_1 ),
    .O(\MASTER/REQ64/$2N3429 )
  );
  X_AND2   \MASTER/REQ64/$2I3431  (
    .I0(\NlwInverterSignal_MASTER/REQ64/$2I3431/I0 ),
    .I1(\MASTER/REQ64/FEEDBACK ),
    .O(\MASTER/REQ64/KO_T_1 )
  );
  X_OR3   \MASTER/REQ64/$2I3411  (
    .I0(\NlwInverterSignal_MASTER/REQ64/$2I3411/I0 ),
    .I1(COMPLETE),
    .I2(\MASTER/REQ64/$2N3399 ),
    .O(\MASTER/REQ64/DONE_0 )
  );
  X_AND2   \MASTER/REQ64/$2I3410  (
    .I0(\MASTER/REQ64/DTO ),
    .I1(NlwRenamedSig_OI_TIME_OUT),
    .O(\MASTER/REQ64/$2N3399 )
  );
  X_OR2   \MASTER/REQ64/$2I3408  (
    .I0(\IIRDY_I- ),
    .I1(\MASTER/IREQ64- ),
    .O(\MASTER/REQ64/INITIAL )
  );
  X_AND2   \MASTER/REQ64/$2I3406  (
    .I0(\NlwInverterSignal_MASTER/REQ64/$2I3406/I0 ),
    .I1(\MASTER/REQ64/FEEDBACK ),
    .O(\MASTER/REQ64/KO_T_0 )
  );
  X_AND2   \MASTER/REQ64/$2I3405  (
    .I0(M_READY),
    .I1(\MASTER/REQ64/$2N3429 ),
    .O(\MASTER/REQ64/$2N3430 )
  );
  X_AND2   \MASTER/REQ64/$2I3394  (
    .I0(\MASTER/REQ64/DTO ),
    .I1(NlwRenamedSig_OI_TIME_OUT),
    .O(\MASTER/REQ64/$2N3396 )
  );
  X_OR3   \MASTER/REQ64/$2I3393  (
    .I0(\NlwInverterSignal_MASTER/REQ64/$2I3393/I0 ),
    .I1(COMPLETE),
    .I2(\MASTER/REQ64/$2N3396 ),
    .O(\MASTER/REQ64/DONE_1 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \MASTER/REQ64/IREQ64-  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(CLK),
    .I(\IREQ64_I- ),
    .O(\MASTER/IREQ64- ),
    .RST(GND)
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \MASTER/REQ64/IREQ64_I-  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(REQ64_CE),
    .CLK(CLK),
    .I(\NS_REQ64- ),
    .O(\IREQ64_I- ),
    .RST(GND)
  );
  X_AND3   \MASTER/REQ64/$1I3616  (
    .I0(\NlwInverterSignal_MASTER/REQ64/$1I3616/I0 ),
    .I1(ADDR_BE),
    .I2(\MASTER/REQUEST64 ),
    .O(\MASTER/REQ64/TURN_ON )
  );
  X_AND2   \MASTER/REQ64/$1I3614  (
    .I0(\NlwInverterSignal_MASTER/REQ64/$1I3614/I0 ),
    .I1(\MASTER/REQ64/FEEDBACK ),
    .O(\MASTER/REQ64/$1N3605 )
  );
  X_AND4   \MASTER/REQ64/$1I3607  (
    .I0(\NlwInverterSignal_MASTER/REQ64/$1I3607/I0 ),
    .I1(\NlwInverterSignal_MASTER/REQ64/$1I3607/I1 ),
    .I2(\NlwInverterSignal_MASTER/REQ64/$1I3607/I2 ),
    .I3(M_DATA_INT),
    .O(\MASTER/REQ64/FEEDBACK )
  );
  X_OR2   \MASTER/REQ64/$1I3569  (
    .I0(\MASTER/REQ64/TURN_ON ),
    .I1(\MASTER/REQ64/$1N3605 ),
    .O(\NlwInverterSignal_MASTER/REQ64/$1I3569/O )
  );
  X_MUX2   \MASTER/REQ64/$1I3568  (
    .IA(\MASTER/REQ64/NS_S_0 ),
    .IB(\MASTER/REQ64/NS_S_1 ),
    .O(\NS_REQ64- ),
    .SEL(STOP_I)
  );
  X_OR2   \MASTER/REQ64/$1I3561  (
    .I0(\MASTER/REQ64/TURN_ON ),
    .I1(\MASTER/REQ64/$1N3615 ),
    .O(\NlwInverterSignal_MASTER/REQ64/$1I3561/O )
  );
  X_AND2   \MASTER/REQ64/$1I3540  (
    .I0(\NlwInverterSignal_MASTER/REQ64/$1I3540/I0 ),
    .I1(ATTEMPT64),
    .O(\MASTER/REQ64/IRDY_64 )
  );
  X_AND4   \MASTER/REQ64/$1I3534  (
    .I0(\NlwInverterSignal_MASTER/REQ64/$1I3534/I0 ),
    .I1(STOP_I),
    .I2(ACK64_I),
    .I3(\MASTER/REQ64/IRDY_64 ),
    .O(\NlwInverterSignal_MASTER/REQ64/$1I3534/O )
  );
  X_BUF   \MASTER/REQ64/$1I3509/NC  (
    .I(\MASTER/REQUEST64 ),
    .O(\NLW_MASTER/REQ64/$1I3509/NC_O_UNCONNECTED )
  );
  X_AND2   \MASTER/REQ64/$1I3562/$1I9  (
    .I0(\MASTER/REQ64/KO_T_1 ),
    .I1(TRDY_M),
    .O(\MASTER/REQ64/$1I3562/M1 )
  );
  X_OR2   \MASTER/REQ64/$1I3562/$1I8  (
    .I0(\MASTER/REQ64/$1I3562/M1 ),
    .I1(\MASTER/REQ64/$1I3562/M0 ),
    .O(\MASTER/REQ64/$1N3615 )
  );
  X_AND2   \MASTER/REQ64/$1I3562/$1I7  (
    .I0(\NlwInverterSignal_MASTER/REQ64/$1I3562/$1I7/I0 ),
    .I1(\MASTER/REQ64/KO_T_0 ),
    .O(\MASTER/REQ64/$1I3562/M0 )
  );
  X_AND2   \MASTER/REQ64/$2I3446/$1I9  (
    .I0(GNT_IN),
    .I1(CFG254),
    .O(\MASTER/REQ64/$2I3446/M1 )
  );
  X_OR2   \MASTER/REQ64/$2I3446/$1I8  (
    .I0(\MASTER/REQ64/$2I3446/M1 ),
    .I1(\MASTER/REQ64/$2I3446/M0 ),
    .O(\MASTER/REQ64/DTO )
  );
  X_AND2   \MASTER/REQ64/$2I3446/$1I7  (
    .I0(\NlwInverterSignal_MASTER/REQ64/$2I3446/$1I7/I0 ),
    .I1(\GNT- ),
    .O(\MASTER/REQ64/$2I3446/M0 )
  );
  X_AND2   \MASTER/XFERFAIL/$1I3027  (
    .I0(FAIL64_INT),
    .I1(M_DATA_INT),
    .O(\MASTER/XFERFAIL/FEEDBACK )
  );
  X_AND3   \MASTER/XFERFAIL/$1I3024  (
    .I0(\NlwInverterSignal_MASTER/XFERFAIL/$1I3024/I0 ),
    .I1(ATTEMPT64),
    .I2(M_DATA_INT),
    .O(\MASTER/XFERFAIL/EQN-X )
  );
  X_AND3   \MASTER/XFERFAIL/$1I3019  (
    .I0(\NlwInverterSignal_MASTER/XFERFAIL/$1I3019/I0 ),
    .I1(ACK64_I),
    .I2(\MASTER/XFERFAIL/EQN-X ),
    .O(\MASTER/XFERFAIL/SET_FAIL64 )
  );
  X_OR2   \MASTER/XFERFAIL/$1I3012  (
    .I0(\MASTER/XFERFAIL/FEEDBACK ),
    .I1(\MASTER/XFERFAIL/SET_FAIL64 ),
    .O(\MASTER/XFERFAIL/NS_0 )
  );
  X_AND2   \MASTER/XFERFAIL/$1I2987  (
    .I0(FAIL64_INT),
    .I1(M_DATA_INT),
    .O(\MASTER/XFERFAIL/NS_1 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \MASTER/XFERFAIL/FAIL_FF  (
    .CE(VCC),
    .CLK(CLK),
    .I(\MASTER/XFERFAIL/NS_FAIL64 ),
    .O(FAIL64_INT),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_MUX2   \MASTER/XFERFAIL/$1I2980  (
    .IA(\MASTER/XFERFAIL/NS_0 ),
    .IB(\MASTER/XFERFAIL/NS_1 ),
    .O(\MASTER/XFERFAIL/NS_FAIL64 ),
    .SEL(TRDY_M)
  );
  X_OR2   \MASTER/OE_FRAME/$8I4093  (
    .I0(\NlwInverterSignal_MASTER/OE_FRAME/$8I4093/I0 ),
    .I1(\MASTER/OE_FRAME/$8N4094 ),
    .O(\MASTER/OE_FRAME/CE_OER )
  );
  X_AND3   \MASTER/OE_FRAME/$8I4089  (
    .I0(\MASTER/REQUEST64 ),
    .I1(SLOT64),
    .I2(ADDR_BE),
    .O(\MASTER/OE_FRAME/$8N4094 )
  );
  X_AND2   \MASTER/OE_FRAME/$8I4077  (
    .I0(\MASTER/REQUEST ),
    .I1(ADDR_BE),
    .O(\MASTER/OE_FRAME/$8N4080 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \MASTER/OE_FRAME/OE_REQ64  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(\MASTER/OE_FRAME/CE_OER ),
    .CLK(CLK),
    .I(\MASTER/OE_FRAME/NS_OER ),
    .O(OE_REQ64),
    .RST(GND)
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \MASTER/OE_FRAME/OE_REQ64_INT  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(\MASTER/OE_FRAME/CE_OER ),
    .CLK(CLK),
    .I(\MASTER/OE_FRAME/NS_OER ),
    .O(\MASTER/OE_FRAME/OE_REQ64_INT_525 ),
    .RST(GND)
  );
  X_MUX2   \MASTER/OE_FRAME/$8I4049  (
    .IA(\MASTER/OE_FRAME/NS_OER_0 ),
    .IB(\MASTER/OE_FRAME/NS_OER_1 ),
    .O(\MASTER/OE_FRAME/NS_OER ),
    .SEL(\MASTER/OE_FRAME/START_AD64 )
  );
  X_OR2   \MASTER/OE_FRAME/$8I4048  (
    .I0(\MASTER/OE_FRAME/MISC64_1 ),
    .I1(\MASTER/OE_FRAME/$8N4025 ),
    .O(\MASTER/OE_FRAME/NS_OER_1 )
  );
  X_AND2   \MASTER/OE_FRAME/$8I4047  (
    .I0(\MASTER/OE_FRAME/MISC64_0 ),
    .I1(\MASTER/OE_FRAME/$8N4018 ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$8I4047/O )
  );
  X_AND2   \MASTER/OE_FRAME/$8I4046  (
    .I0(\MASTER/OE_FRAME/$8N4024 ),
    .I1(\IREQ64_I- ),
    .O(\MASTER/OE_FRAME/$8N4025 )
  );
  X_OR2   \MASTER/OE_FRAME/$8I4045  (
    .I0(\NlwInverterSignal_MASTER/OE_FRAME/$8I4045/I0 ),
    .I1(\NlwInverterSignal_MASTER/OE_FRAME/$8I4045/I1 ),
    .O(\MASTER/OE_FRAME/$8N4024 )
  );
  X_OR2   \MASTER/OE_FRAME/$8I4044  (
    .I0(\NlwInverterSignal_MASTER/OE_FRAME/$8I4044/I0 ),
    .I1(\NlwInverterSignal_MASTER/OE_FRAME/$8I4044/I1 ),
    .O(\MASTER/OE_FRAME/$8N4019 )
  );
  X_AND2   \MASTER/OE_FRAME/$8I4043  (
    .I0(\MASTER/OE_FRAME/$8N4019 ),
    .I1(\IREQ64_I- ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$8I4043/O )
  );
  X_OR2   \MASTER/OE_FRAME/$8I4007  (
    .I0(\NlwInverterSignal_MASTER/OE_FRAME/$8I4007/I0 ),
    .I1(\MASTER/OE_FRAME/$8N4080 ),
    .O(\MASTER/OE_FRAME/CE_OEF )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \MASTER/OE_FRAME/OE_FRAME_INT  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(\MASTER/OE_FRAME/CE_OEF ),
    .CLK(CLK),
    .I(\MASTER/OE_FRAME/NS_OEF ),
    .O(\MASTER/OE_FRAME/OE_FRAME_INT_509 ),
    .RST(GND)
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \MASTER/OE_FRAME/OE_FRAME  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(\MASTER/OE_FRAME/CE_OEF ),
    .CLK(CLK),
    .I(\MASTER/OE_FRAME/NS_OEF ),
    .O(OE_FRAME),
    .RST(GND)
  );
  X_AND2   \MASTER/OE_FRAME/$8I3975  (
    .I0(\MASTER/OE_FRAME/$8N3991 ),
    .I1(\IFRAME_I- ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$8I3975/O )
  );
  X_OR2   \MASTER/OE_FRAME/$8I3974  (
    .I0(\NlwInverterSignal_MASTER/OE_FRAME/$8I3974/I0 ),
    .I1(\NlwInverterSignal_MASTER/OE_FRAME/$8I3974/I1 ),
    .O(\MASTER/OE_FRAME/$8N3991 )
  );
  X_OR2   \MASTER/OE_FRAME/$8I3973  (
    .I0(\NlwInverterSignal_MASTER/OE_FRAME/$8I3973/I0 ),
    .I1(\NlwInverterSignal_MASTER/OE_FRAME/$8I3973/I1 ),
    .O(\MASTER/OE_FRAME/$8N3986 )
  );
  X_AND2   \MASTER/OE_FRAME/$8I3972  (
    .I0(\MASTER/OE_FRAME/$8N3986 ),
    .I1(\IFRAME_I- ),
    .O(\MASTER/OE_FRAME/$8N3985 )
  );
  X_AND2   \MASTER/OE_FRAME/$8I3971  (
    .I0(\MASTER/OE_FRAME/MISC_0 ),
    .I1(\MASTER/OE_FRAME/$8N3992 ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$8I3971/O )
  );
  X_OR2   \MASTER/OE_FRAME/$8I3970  (
    .I0(\MASTER/OE_FRAME/MISC_1 ),
    .I1(\MASTER/OE_FRAME/$8N3985 ),
    .O(\MASTER/OE_FRAME/NS_OEF_1 )
  );
  X_MUX2   \MASTER/OE_FRAME/$8I3969  (
    .IA(\MASTER/OE_FRAME/NS_OEF_0 ),
    .IB(\MASTER/OE_FRAME/NS_OEF_1 ),
    .O(\MASTER/OE_FRAME/NS_OEF ),
    .SEL(\MASTER/OE_FRAME/START_AD )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \MASTER/OE_FRAME/OE_IRDY  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(CLK),
    .I(\MASTER/OE_FRAME/OE_FRAME_INT_509 ),
    .O(OE_IRDY),
    .RST(GND)
  );
  X_MUX2   \MASTER/OE_FRAME/$7I3978  (
    .IA(\MASTER/OE_FRAME/NS64_0 ),
    .IB(\MASTER/OE_FRAME/NS64_1 ),
    .O(\MASTER/OE_FRAME/NS64 ),
    .SEL(\MASTER/OE_FRAME/START_AD64 )
  );
  X_OR2   \MASTER/OE_FRAME/$7I3977  (
    .I0(\MASTER/OE_FRAME/MISC64_1 ),
    .I1(\MASTER/OE_FRAME/$7N3953 ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$7I3977/O )
  );
  X_AND2   \MASTER/OE_FRAME/$7I3976  (
    .I0(\IREQ64_I- ),
    .I1(\MASTER/DEV_TO ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$7I3976/O )
  );
  X_OR2   \MASTER/OE_FRAME/$7I3975  (
    .I0(\NlwInverterSignal_MASTER/OE_FRAME/$7I3975/I0 ),
    .I1(\NlwInverterSignal_MASTER/OE_FRAME/$7I3975/I1 ),
    .O(\MASTER/OE_FRAME/$7N3955 )
  );
  X_AND2   \MASTER/OE_FRAME/$7I3974  (
    .I0(\MASTER/OE_FRAME/MISC64_0 ),
    .I1(\MASTER/OE_FRAME/$7N3936 ),
    .O(\MASTER/OE_FRAME/NS64_0 )
  );
  X_AND2   \MASTER/OE_FRAME/$7I3973  (
    .I0(\MASTER/OE_FRAME/$7N3948 ),
    .I1(\IREQ64_I- ),
    .O(\MASTER/OE_FRAME/$7N3953 )
  );
  X_AND2   \MASTER/OE_FRAME/$7I3972  (
    .I0(\IREQ64_I- ),
    .I1(\MASTER/DEV_TO ),
    .O(\MASTER/OE_FRAME/MISC64_3 )
  );
  X_OR2   \MASTER/OE_FRAME/$7I3971  (
    .I0(\MASTER/OE_FRAME/$7N3952 ),
    .I1(\MASTER/OE_FRAME/MISC64_3 ),
    .O(\MASTER/OE_FRAME/MISC64_1 )
  );
  X_AND2   \MASTER/OE_FRAME/$7I3970  (
    .I0(\MASTER/OE_FRAME/OE_REQ64_INT_525 ),
    .I1(GNT_IN),
    .O(\MASTER/OE_FRAME/$7N3947 )
  );
  X_AND2   \MASTER/OE_FRAME/$7I3969  (
    .I0(GNT_IN),
    .I1(\MASTER/OE_FRAME/DR_BUS1 ),
    .O(\MASTER/OE_FRAME/$7N3949 )
  );
  X_OR2   \MASTER/OE_FRAME/$7I3968  (
    .I0(\NlwInverterSignal_MASTER/OE_FRAME/$7I3968/I0 ),
    .I1(\NlwInverterSignal_MASTER/OE_FRAME/$7I3968/I1 ),
    .O(\MASTER/OE_FRAME/$7N3948 )
  );
  X_OR2   \MASTER/OE_FRAME/$7I3967  (
    .I0(\MASTER/OE_FRAME/$7N3949 ),
    .I1(\MASTER/OE_FRAME/$7N3947 ),
    .O(\MASTER/OE_FRAME/$7N3952 )
  );
  X_OR2   \MASTER/OE_FRAME/$7I3966  (
    .I0(\NlwInverterSignal_MASTER/OE_FRAME/$7I3966/I0 ),
    .I1(\NlwInverterSignal_MASTER/OE_FRAME/$7I3966/I1 ),
    .O(\MASTER/OE_FRAME/$7N3940 )
  );
  X_AND2   \MASTER/OE_FRAME/$7I3965  (
    .I0(\MASTER/OE_FRAME/$7N3940 ),
    .I1(\IREQ64_I- ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$7I3965/O )
  );
  X_AND3   \MASTER/OE_FRAME/$7I3964  (
    .I0(\MASTER/OE_FRAME/SLOT64 ),
    .I1(\MASTER/OE_FRAME/$7N3955 ),
    .I2(\MASTER/OE_FRAME/MISC64_2 ),
    .O(\MASTER/OE_FRAME/MISC64_0 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \MASTER/OE_FRAME/SLOT64_FF  (
    .CE(VCC),
    .CLK(CLK),
    .I(\MASTER/OE_FRAME/NS64 ),
    .O(\MASTER/OE_FRAME/SLOT64 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_MUX2   \MASTER/OE_FRAME/$6I3741  (
    .IA(\MASTER/OE_FRAME/NS_0 ),
    .IB(\MASTER/OE_FRAME/NS_1 ),
    .O(\MASTER/OE_FRAME/NS ),
    .SEL(\MASTER/OE_FRAME/START_AD )
  );
  X_OR2   \MASTER/OE_FRAME/$6I3740  (
    .I0(\MASTER/OE_FRAME/MISC_1 ),
    .I1(\MASTER/OE_FRAME/$6N3723 ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$6I3740/O )
  );
  X_AND2   \MASTER/OE_FRAME/$6I3739  (
    .I0(\IFRAME_I- ),
    .I1(\MASTER/DEV_TO ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$6I3739/O )
  );
  X_OR2   \MASTER/OE_FRAME/$6I3738  (
    .I0(\NlwInverterSignal_MASTER/OE_FRAME/$6I3738/I0 ),
    .I1(\NlwInverterSignal_MASTER/OE_FRAME/$6I3738/I1 ),
    .O(\MASTER/OE_FRAME/$6N3725 )
  );
  X_AND2   \MASTER/OE_FRAME/$6I3737  (
    .I0(\MASTER/OE_FRAME/MISC_0 ),
    .I1(\MASTER/OE_FRAME/$6N3707 ),
    .O(\MASTER/OE_FRAME/NS_0 )
  );
  X_AND2   \MASTER/OE_FRAME/$6I3736  (
    .I0(\MASTER/OE_FRAME/$6N3718 ),
    .I1(\IFRAME_I- ),
    .O(\MASTER/OE_FRAME/$6N3723 )
  );
  X_AND2   \MASTER/OE_FRAME/$6I3735  (
    .I0(\IFRAME_I- ),
    .I1(\MASTER/DEV_TO ),
    .O(\MASTER/OE_FRAME/MISC_3 )
  );
  X_OR2   \MASTER/OE_FRAME/$6I3734  (
    .I0(\MASTER/OE_FRAME/$6N3722 ),
    .I1(\MASTER/OE_FRAME/MISC_3 ),
    .O(\MASTER/OE_FRAME/MISC_1 )
  );
  X_AND2   \MASTER/OE_FRAME/$6I3733  (
    .I0(\MASTER/OE_FRAME/OE_FRAME_INT_509 ),
    .I1(GNT_IN),
    .O(\MASTER/OE_FRAME/$6N3717 )
  );
  X_AND2   \MASTER/OE_FRAME/$6I3732  (
    .I0(GNT_IN),
    .I1(\MASTER/OE_FRAME/DR_BUS1 ),
    .O(\MASTER/OE_FRAME/$6N3719 )
  );
  X_OR2   \MASTER/OE_FRAME/$6I3731  (
    .I0(\NlwInverterSignal_MASTER/OE_FRAME/$6I3731/I0 ),
    .I1(\NlwInverterSignal_MASTER/OE_FRAME/$6I3731/I1 ),
    .O(\MASTER/OE_FRAME/$6N3718 )
  );
  X_OR2   \MASTER/OE_FRAME/$6I3730  (
    .I0(\MASTER/OE_FRAME/$6N3719 ),
    .I1(\MASTER/OE_FRAME/$6N3717 ),
    .O(\MASTER/OE_FRAME/$6N3722 )
  );
  X_OR2   \MASTER/OE_FRAME/$6I3729  (
    .I0(\NlwInverterSignal_MASTER/OE_FRAME/$6I3729/I0 ),
    .I1(\NlwInverterSignal_MASTER/OE_FRAME/$6I3729/I1 ),
    .O(\MASTER/OE_FRAME/$6N3710 )
  );
  X_AND2   \MASTER/OE_FRAME/$6I3728  (
    .I0(\MASTER/OE_FRAME/$6N3710 ),
    .I1(\IFRAME_I- ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$6I3728/O )
  );
  X_AND3   \MASTER/OE_FRAME/$6I3727  (
    .I0(\MASTER/OE_FRAME/SLOT ),
    .I1(\MASTER/OE_FRAME/$6N3725 ),
    .I2(\MASTER/OE_FRAME/MISC_2 ),
    .O(\MASTER/OE_FRAME/MISC_0 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \MASTER/OE_FRAME/SLOT_FF  (
    .CE(VCC),
    .CLK(CLK),
    .I(\MASTER/OE_FRAME/NS ),
    .O(\MASTER/OE_FRAME/SLOT ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \MASTER/OE_FRAME/H_PAR_OE  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(CLK),
    .I(NlwRenamedSig_OI_OE_ADO_B64),
    .O(NlwRenamedSig_OI_OE_PAR64),
    .RST(GND)
  );
  X_OR2   \MASTER/OE_FRAME/$5I3899  (
    .I0(\NlwInverterSignal_MASTER/OE_FRAME/$5I3899/I0 ),
    .I1(\MASTER/OE_FRAME/$5N3870 ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$5I3899/O )
  );
  X_AND2   \MASTER/OE_FRAME/$5I3898  (
    .I0(\NlwInverterSignal_MASTER/OE_FRAME/$5I3898/I0 ),
    .I1(\NlwInverterSignal_MASTER/OE_FRAME/$5I3898/I1 ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$5I3898/O )
  );
  X_OR2   \MASTER/OE_FRAME/$5I3893  (
    .I0(\NlwInverterSignal_MASTER/OE_FRAME/$5I3893/I0 ),
    .I1(\MASTER/OE_FRAME/START_AD64 ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$5I3893/O )
  );
  X_AND2   \MASTER/OE_FRAME/$5I3891  (
    .I0(\NlwInverterSignal_MASTER/OE_FRAME/$5I3891/I0 ),
    .I1(\MASTER/OE_FRAME/SLOT64 ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$5I3891/O )
  );
  X_OR2   \MASTER/OE_FRAME/$5I3890  (
    .I0(\NlwInverterSignal_MASTER/OE_FRAME/$5I3890/I0 ),
    .I1(\MASTER/OE_FRAME/START_AD64 ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$5I3890/O )
  );
  X_OR2   \MASTER/OE_FRAME/$5I3889  (
    .I0(\NlwInverterSignal_MASTER/OE_FRAME/$5I3889/I0 ),
    .I1(\MASTER/OE_FRAME/START_AD64 ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$5I3889/O )
  );
  X_OR2   \MASTER/OE_FRAME/$5I3888  (
    .I0(\NlwInverterSignal_MASTER/OE_FRAME/$5I3888/I0 ),
    .I1(\MASTER/OE_FRAME/START_AD64 ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$5I3888/O )
  );
  X_OR2   \MASTER/OE_FRAME/$5I3887  (
    .I0(\NlwInverterSignal_MASTER/OE_FRAME/$5I3887/I0 ),
    .I1(\MASTER/OE_FRAME/START_AD64 ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$5I3887/O )
  );
  X_OR2   \MASTER/OE_FRAME/$5I3886  (
    .I0(\NlwInverterSignal_MASTER/OE_FRAME/$5I3886/I0 ),
    .I1(\MASTER/OE_FRAME/$5N3869 ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$5I3886/O )
  );
  X_OR2   \MASTER/OE_FRAME/$5I3885  (
    .I0(\NlwInverterSignal_MASTER/OE_FRAME/$5I3885/I0 ),
    .I1(\MASTER/OE_FRAME/$5N3868 ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$5I3885/O )
  );
  X_OR2   \MASTER/OE_FRAME/$5I3884  (
    .I0(\NlwInverterSignal_MASTER/OE_FRAME/$5I3884/I0 ),
    .I1(\MASTER/OE_FRAME/$5N3874 ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$5I3884/O )
  );
  X_AND2   \MASTER/OE_FRAME/$5I3883  (
    .I0(\NlwInverterSignal_MASTER/OE_FRAME/$5I3883/I0 ),
    .I1(\NlwInverterSignal_MASTER/OE_FRAME/$5I3883/I1 ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$5I3883/O )
  );
  X_AND2   \MASTER/OE_FRAME/$5I3882  (
    .I0(\NlwInverterSignal_MASTER/OE_FRAME/$5I3882/I0 ),
    .I1(\NlwInverterSignal_MASTER/OE_FRAME/$5I3882/I1 ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$5I3882/O )
  );
  X_AND2   \MASTER/OE_FRAME/$5I3881  (
    .I0(\NlwInverterSignal_MASTER/OE_FRAME/$5I3881/I0 ),
    .I1(\NlwInverterSignal_MASTER/OE_FRAME/$5I3881/I1 ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$5I3881/O )
  );
  X_AND2   \MASTER/OE_FRAME/$5I3880  (
    .I0(M_WRDN),
    .I1(\MASTER/OE_FRAME/SLOT64 ),
    .O(\MASTER/OE_FRAME/$5N3874 )
  );
  X_AND2   \MASTER/OE_FRAME/$5I3879  (
    .I0(M_WRDN),
    .I1(\MASTER/OE_FRAME/SLOT64 ),
    .O(\MASTER/OE_FRAME/$5N3869 )
  );
  X_AND2   \MASTER/OE_FRAME/$5I3878  (
    .I0(M_WRDN),
    .I1(\MASTER/OE_FRAME/SLOT64 ),
    .O(\MASTER/OE_FRAME/$5N3868 )
  );
  X_AND2   \MASTER/OE_FRAME/$5I3877  (
    .I0(M_WRDN),
    .I1(\MASTER/OE_FRAME/SLOT64 ),
    .O(\MASTER/OE_FRAME/$5N3870 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \MASTER/OE_FRAME/L_PAR_OE  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(CLK),
    .I(NlwRenamedSig_OI_OE_ADO_B),
    .O(NlwRenamedSig_OI_OE_PAR),
    .RST(GND)
  );
  X_AND2   \MASTER/OE_FRAME/$4I3785  (
    .I0(\NlwInverterSignal_MASTER/OE_FRAME/$4I3785/I0 ),
    .I1(\MASTER/OE_FRAME/SLOT ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$4I3785/O )
  );
  X_OR2   \MASTER/OE_FRAME/$4I3784  (
    .I0(\NlwInverterSignal_MASTER/OE_FRAME/$4I3784/I0 ),
    .I1(\MASTER/OE_FRAME/START_AD ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$4I3784/O )
  );
  X_OR2   \MASTER/OE_FRAME/$4I3783  (
    .I0(\NlwInverterSignal_MASTER/OE_FRAME/$4I3783/I0 ),
    .I1(\MASTER/OE_FRAME/START_AD ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$4I3783/O )
  );
  X_OR2   \MASTER/OE_FRAME/$4I3782  (
    .I0(\NlwInverterSignal_MASTER/OE_FRAME/$4I3782/I0 ),
    .I1(\MASTER/OE_FRAME/START_AD ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$4I3782/O )
  );
  X_OR2   \MASTER/OE_FRAME/$4I3781  (
    .I0(\NlwInverterSignal_MASTER/OE_FRAME/$4I3781/I0 ),
    .I1(\MASTER/OE_FRAME/START_AD ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$4I3781/O )
  );
  X_OR2   \MASTER/OE_FRAME/$4I3780  (
    .I0(\NlwInverterSignal_MASTER/OE_FRAME/$4I3780/I0 ),
    .I1(\MASTER/OE_FRAME/START_AD ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$4I3780/O )
  );
  X_AND2   \MASTER/OE_FRAME/$4I3779  (
    .I0(\NlwInverterSignal_MASTER/OE_FRAME/$4I3779/I0 ),
    .I1(\NlwInverterSignal_MASTER/OE_FRAME/$4I3779/I1 ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$4I3779/O )
  );
  X_OR2   \MASTER/OE_FRAME/$4I3778  (
    .I0(\NlwInverterSignal_MASTER/OE_FRAME/$4I3778/I0 ),
    .I1(\MASTER/OE_FRAME/$4N3740 ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$4I3778/O )
  );
  X_OR2   \MASTER/OE_FRAME/$4I3776  (
    .I0(\NlwInverterSignal_MASTER/OE_FRAME/$4I3776/I0 ),
    .I1(\MASTER/OE_FRAME/$4N3739 ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$4I3776/O )
  );
  X_OR2   \MASTER/OE_FRAME/$4I3774  (
    .I0(\NlwInverterSignal_MASTER/OE_FRAME/$4I3774/I0 ),
    .I1(\MASTER/OE_FRAME/$4N3738 ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$4I3774/O )
  );
  X_OR2   \MASTER/OE_FRAME/$4I3772  (
    .I0(\NlwInverterSignal_MASTER/OE_FRAME/$4I3772/I0 ),
    .I1(\MASTER/OE_FRAME/$4N3749 ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$4I3772/O )
  );
  X_AND2   \MASTER/OE_FRAME/$4I3770  (
    .I0(\NlwInverterSignal_MASTER/OE_FRAME/$4I3770/I0 ),
    .I1(\NlwInverterSignal_MASTER/OE_FRAME/$4I3770/I1 ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$4I3770/O )
  );
  X_AND2   \MASTER/OE_FRAME/$4I3769  (
    .I0(\NlwInverterSignal_MASTER/OE_FRAME/$4I3769/I0 ),
    .I1(\NlwInverterSignal_MASTER/OE_FRAME/$4I3769/I1 ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$4I3769/O )
  );
  X_AND2   \MASTER/OE_FRAME/$4I3768  (
    .I0(\NlwInverterSignal_MASTER/OE_FRAME/$4I3768/I0 ),
    .I1(\NlwInverterSignal_MASTER/OE_FRAME/$4I3768/I1 ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$4I3768/O )
  );
  X_AND2   \MASTER/OE_FRAME/$4I3767  (
    .I0(M_WRDN),
    .I1(\MASTER/OE_FRAME/SLOT ),
    .O(\MASTER/OE_FRAME/$4N3749 )
  );
  X_AND2   \MASTER/OE_FRAME/$4I3766  (
    .I0(M_WRDN),
    .I1(\MASTER/OE_FRAME/SLOT ),
    .O(\MASTER/OE_FRAME/$4N3739 )
  );
  X_AND2   \MASTER/OE_FRAME/$4I3765  (
    .I0(M_WRDN),
    .I1(\MASTER/OE_FRAME/SLOT ),
    .O(\MASTER/OE_FRAME/$4N3738 )
  );
  X_AND2   \MASTER/OE_FRAME/$4I3764  (
    .I0(M_WRDN),
    .I1(\MASTER/OE_FRAME/SLOT ),
    .O(\MASTER/OE_FRAME/$4N3740 )
  );
  X_AND2   \MASTER/OE_FRAME/$3I3110  (
    .I0(PERR_EN),
    .I1(M_DATA_INT),
    .O(\MASTER/OE_FRAME/EQN-A )
  );
  X_AND4   \MASTER/OE_FRAME/$3I3105  (
    .I0(\NlwInverterSignal_MASTER/OE_FRAME/$3I3105/I0 ),
    .I1(\NlwInverterSignal_MASTER/OE_FRAME/$3I3105/I1 ),
    .I2(\NlwInverterSignal_MASTER/OE_FRAME/$3I3105/I2 ),
    .I3(\MASTER/OE_FRAME/EQN-A ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$3I3105/O )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \MASTER/OE_FRAME/I_PERR_HOLD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(CLK),
    .I(\MASTER/OE_FRAME/SET_OE_PERR ),
    .O(\MASTER/OE_FRAME/HOLD_OE_PERR ),
    .RST(GND)
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \MASTER/OE_FRAME/PERR_OE  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(CLK),
    .I(\MASTER/OE_FRAME/NS_OE_PERR ),
    .O(OE_PERR),
    .RST(GND)
  );
  X_OR3   \MASTER/OE_FRAME/$3I3093  (
    .I0(\NlwInverterSignal_MASTER/OE_FRAME/$3I3093/I0 ),
    .I1(\NlwInverterSignal_MASTER/OE_FRAME/$3I3093/I1 ),
    .I2(\NlwInverterSignal_MASTER/OE_FRAME/$3I3093/I2 ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$3I3093/O )
  );
  X_AND4   \MASTER/OE_FRAME/$2I3723  (
    .I0(\NlwInverterSignal_MASTER/OE_FRAME/$2I3723/I0 ),
    .I1(\FRAME- ),
    .I2(\IRDY- ),
    .I3(\MASTER/OE_FRAME/REQUEST64Q ),
    .O(\MASTER/OE_FRAME/START_AD64 )
  );
  X_AND4   \MASTER/OE_FRAME/$2I3711  (
    .I0(\NlwInverterSignal_MASTER/OE_FRAME/$2I3711/I0 ),
    .I1(\FRAME- ),
    .I2(\IRDY- ),
    .I3(\MASTER/OE_FRAME/REQUESTQ ),
    .O(\MASTER/OE_FRAME/START_AD )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \MASTER/OE_FRAME/$1I3713  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(CLK),
    .I(\MASTER/OE_FRAME/$1N3716 ),
    .O(\MASTER/OE_FRAME/DUMMY ),
    .RST(GND)
  );
  X_INV   \MASTER/OE_FRAME/$1I3701  (
    .I(\$1N4834 ),
    .O(\MASTER/OE_FRAME/$1N3703 )
  );
  X_OR3   \MASTER/OE_FRAME/$1I3697  (
    .I0(DR_BUS_INT),
    .I1(\MASTER/OE_FRAME/DR_BUSQ ),
    .I2(\MASTER/OE_FRAME/DUMMY ),
    .O(\MASTER/OE_FRAME/DR_BUS1 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \MASTER/OE_FRAME/$1I3695  (
    .CE(\MASTER/OE_FRAME/$1N3703 ),
    .CLK(CLK),
    .I(DR_BUS_INT),
    .O(\MASTER/OE_FRAME/DR_BUSQ ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \MASTER/OE_FRAME/$1I3693  (
    .CE(VCC),
    .CLK(CLK),
    .I(\MASTER/REQUEST64 ),
    .O(\MASTER/OE_FRAME/REQUEST64Q ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \MASTER/OE_FRAME/$1I3692  (
    .CE(VCC),
    .CLK(CLK),
    .I(\MASTER/OE_FRAME/$1N3685 ),
    .O(\MASTER/OE_FRAME/REQUESTQ ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_ONE   \MASTER/OE_FRAME/$1I3691/$1I2220  (
    .O(\MASTER/OE_FRAME/$1I3691/$1N2216 )
  );
  X_BUF   \MASTER/OE_FRAME/$1I3691/H  (
    .I(\MASTER/OE_FRAME/$1I3691/$1N2216 ),
    .O(\MASTER/OE_FRAME/$1N3685 )
  );
  X_ZERO   \MASTER/OE_FRAME/$1I3717/$1I2218  (
    .O(\MASTER/OE_FRAME/$1I3717/$1N2216 )
  );
  X_BUF   \MASTER/OE_FRAME/$1I3717/L  (
    .I(\MASTER/OE_FRAME/$1I3717/$1N2216 ),
    .O(\MASTER/OE_FRAME/$1N3716 )
  );
  X_AND2   \MASTER/OE_FRAME/$5I4044/$1I9  (
    .I0(\MASTER/OE_FRAME/$5N3892 ),
    .I1(SLOT64),
    .O(\MASTER/OE_FRAME/$5I4044/M1 )
  );
  X_OR2   \MASTER/OE_FRAME/$5I4044/$1I8  (
    .I0(\MASTER/OE_FRAME/$5I4044/M1 ),
    .I1(\MASTER/OE_FRAME/$5I4044/M0 ),
    .O(NlwRenamedSig_OI_OE_ADO_T64)
  );
  X_AND2   \MASTER/OE_FRAME/$5I4044/$1I7  (
    .I0(\NlwInverterSignal_MASTER/OE_FRAME/$5I4044/$1I7/I0 ),
    .I1(\NlwInverterSignal_MASTER/OE_FRAME/$5I4044/$1I7/I1 ),
    .O(\MASTER/OE_FRAME/$5I4044/M0 )
  );
  X_AND2   \MASTER/OE_FRAME/$5I4045/$1I9  (
    .I0(\MASTER/OE_FRAME/$5N3873 ),
    .I1(SLOT64),
    .O(\MASTER/OE_FRAME/$5I4045/M1 )
  );
  X_OR2   \MASTER/OE_FRAME/$5I4045/$1I8  (
    .I0(\MASTER/OE_FRAME/$5I4045/M1 ),
    .I1(\MASTER/OE_FRAME/$5I4045/M0 ),
    .O(NlwRenamedSig_OI_OE_ADO_LT64)
  );
  X_AND2   \MASTER/OE_FRAME/$5I4045/$1I7  (
    .I0(\NlwInverterSignal_MASTER/OE_FRAME/$5I4045/$1I7/I0 ),
    .I1(\NlwInverterSignal_MASTER/OE_FRAME/$5I4045/$1I7/I1 ),
    .O(\MASTER/OE_FRAME/$5I4045/M0 )
  );
  X_AND2   \MASTER/OE_FRAME/$5I4046/$1I9  (
    .I0(\MASTER/OE_FRAME/$5N3872 ),
    .I1(SLOT64),
    .O(\MASTER/OE_FRAME/$5I4046/M1 )
  );
  X_OR2   \MASTER/OE_FRAME/$5I4046/$1I8  (
    .I0(\MASTER/OE_FRAME/$5I4046/M1 ),
    .I1(\MASTER/OE_FRAME/$5I4046/M0 ),
    .O(NlwRenamedSig_OI_OE_ADO_LB64)
  );
  X_AND2   \MASTER/OE_FRAME/$5I4046/$1I7  (
    .I0(\NlwInverterSignal_MASTER/OE_FRAME/$5I4046/$1I7/I0 ),
    .I1(\NlwInverterSignal_MASTER/OE_FRAME/$5I4046/$1I7/I1 ),
    .O(\MASTER/OE_FRAME/$5I4046/M0 )
  );
  X_AND2   \MASTER/OE_FRAME/$5I4047/$1I9  (
    .I0(\MASTER/OE_FRAME/$5N3871 ),
    .I1(SLOT64),
    .O(\MASTER/OE_FRAME/$5I4047/M1 )
  );
  X_OR2   \MASTER/OE_FRAME/$5I4047/$1I8  (
    .I0(\MASTER/OE_FRAME/$5I4047/M1 ),
    .I1(\MASTER/OE_FRAME/$5I4047/M0 ),
    .O(NlwRenamedSig_OI_OE_ADO_B64)
  );
  X_AND2   \MASTER/OE_FRAME/$5I4047/$1I7  (
    .I0(\NlwInverterSignal_MASTER/OE_FRAME/$5I4047/$1I7/I0 ),
    .I1(\NlwInverterSignal_MASTER/OE_FRAME/$5I4047/$1I7/I1 ),
    .O(\MASTER/OE_FRAME/$5I4047/M0 )
  );
  X_AND2   \MASTER/OE_FRAME/$5I4048/$1I9  (
    .I0(\MASTER/OE_FRAME/$5N3876 ),
    .I1(SLOT64),
    .O(\MASTER/OE_FRAME/$5I4048/M1 )
  );
  X_OR2   \MASTER/OE_FRAME/$5I4048/$1I8  (
    .I0(\MASTER/OE_FRAME/$5I4048/M1 ),
    .I1(\MASTER/OE_FRAME/$5I4048/M0 ),
    .O(NlwRenamedSig_OI_OE_CBE64)
  );
  X_AND2   \MASTER/OE_FRAME/$5I4048/$1I7  (
    .I0(\NlwInverterSignal_MASTER/OE_FRAME/$5I4048/$1I7/I0 ),
    .I1(\NlwInverterSignal_MASTER/OE_FRAME/$5I4048/$1I7/I1 ),
    .O(\MASTER/OE_FRAME/$5I4048/M0 )
  );
  X_OR2   \MASTER/S_TAR/$1I2605  (
    .I0(\NlwInverterSignal_MASTER/S_TAR/$1I2605/I0 ),
    .I1(\MASTER/DEV_TO ),
    .O(\MASTER/S_TAR/$1N2602 )
  );
  X_AND3   \MASTER/S_TAR/$1I2601  (
    .I0(\IFRAME_I- ),
    .I1(M_DATA_INT),
    .I2(\MASTER/S_TAR/$1N2602 ),
    .O(\MASTER/S_TAR/NS_S_TAR )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \MASTER/S_TAR/S_TAR  (
    .CE(VCC),
    .CLK(CLK),
    .I(\MASTER/S_TAR/NS_S_TAR ),
    .O(\MASTER/S_TAR ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_INV   \MASTER/DEV_TO/$1I2836  (
    .I(M_DATA_INT),
    .O(\MASTER/DEV_TO/$1N2840 )
  );
  X_AND2   \MASTER/DEV_TO/$1I2833  (
    .I0(\MASTER/DEV_TO/WAS_NO_RESPONSE ),
    .I1(\MASTER/DEV_TO/WAS_SUBTRACTIVE ),
    .O(\MASTER/DEV_TO )
  );
  X_AND2   \MASTER/DEV_TO/$1I2823  (
    .I0(\DEVSEL- ),
    .I1(\MASTER/DEV_TO/PASS_TO ),
    .O(\MASTER/DEV_TO/WAS_NO_RESPONSE )
  );
  X_INV   \MASTER/DEV_TO/$1I2819  (
    .I(\DEVSEL- ),
    .O(\MASTER/DEV_TO/$1N2820 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \MASTER/DEV_TO/$1I2807  (
    .CE(VCC),
    .CLK(CLK),
    .I(\MASTER/DEV_TO/WAS_MEDIUM ),
    .O(\MASTER/DEV_TO/WAS_SLOW ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \MASTER/DEV_TO/$1I2803  (
    .CE(VCC),
    .CLK(CLK),
    .I(\MASTER/DEV_TO/WAS_FAST ),
    .O(\MASTER/DEV_TO/WAS_MEDIUM ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \MASTER/DEV_TO/$1I2799  (
    .CE(VCC),
    .CLK(CLK),
    .I(\MASTER/DEV_TO/FAST ),
    .O(\MASTER/DEV_TO/WAS_FAST ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \MASTER/DEV_TO/$1I2796  (
    .CE(VCC),
    .CLK(CLK),
    .I(\MASTER/DEV_TO/ADDR ),
    .O(\MASTER/DEV_TO/FAST ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND2   \MASTER/DEV_TO/$1I2789  (
    .I0(\NlwInverterSignal_MASTER/DEV_TO/$1I2789/I0 ),
    .I1(\MASTER/IFRAME- ),
    .O(\MASTER/DEV_TO/ADDR )
  );
  X_OR2   \MASTER/DEV_TO/$1I2816/$1I2214  (
    .I0(\MASTER/DEV_TO/ADDR ),
    .I1(\MASTER/DEV_TO/PASS_TO ),
    .O(\MASTER/DEV_TO/$1I2816/$1N2215 )
  );
  X_AND2   \MASTER/DEV_TO/$1I2816/$1I2213  (
    .I0(\NlwInverterSignal_MASTER/DEV_TO/$1I2816/$1I2213/I0 ),
    .I1(\MASTER/DEV_TO/$1I2816/$1N2215 ),
    .O(\MASTER/DEV_TO/$1I2816/D )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \MASTER/DEV_TO/$1I2816/FDCE  (
    .CE(VCC),
    .CLK(CLK),
    .I(\MASTER/DEV_TO/$1I2816/D ),
    .O(\MASTER/DEV_TO/PASS_TO ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_OR2   \MASTER/DEV_TO/$1I2838/$1I2214  (
    .I0(\MASTER/DEV_TO/WAS_SLOW ),
    .I1(\MASTER/DEV_TO/WAS_SUBTRACTIVE ),
    .O(\MASTER/DEV_TO/$1I2838/$1N2215 )
  );
  X_AND2   \MASTER/DEV_TO/$1I2838/$1I2213  (
    .I0(\NlwInverterSignal_MASTER/DEV_TO/$1I2838/$1I2213/I0 ),
    .I1(\MASTER/DEV_TO/$1I2838/$1N2215 ),
    .O(\MASTER/DEV_TO/$1I2838/D )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \MASTER/DEV_TO/$1I2838/FDCE  (
    .CE(VCC),
    .CLK(CLK),
    .I(\MASTER/DEV_TO/$1I2838/D ),
    .O(\MASTER/DEV_TO/WAS_SUBTRACTIVE ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_INV   \MASTER/$4I3071/INV1  (
    .I(M_CBE1),
    .O(\MASTER/$4I3071/$1N2280 )
  );
  X_INV   \MASTER/$4I3071/INV2  (
    .I(M_CBE2),
    .O(\MASTER/$4I3071/$1N2278 )
  );
  X_INV   \MASTER/$4I3071/INV3  (
    .I(M_CBE3),
    .O(\MASTER/$4I3071/$1N2277 )
  );
  X_AND4   \MASTER/$4I3071/AND4  (
    .I0(M_CBE0),
    .I1(\MASTER/$4I3071/$1N2280 ),
    .I2(\MASTER/$4I3071/$1N2278 ),
    .I3(\MASTER/$4I3071/$1N2277 ),
    .O(\MASTER/$4N3021 )
  );
  X_BUF   \MASTER/$4I3125/NC  (
    .I(M_CBE7),
    .O(\NLW_MASTER/$4I3125/NC_O_UNCONNECTED )
  );
  X_BUF   \MASTER/$4I3126/NC  (
    .I(M_CBE6),
    .O(\NLW_MASTER/$4I3126/NC_O_UNCONNECTED )
  );
  X_BUF   \MASTER/$4I3127/NC  (
    .I(M_CBE5),
    .O(\NLW_MASTER/$4I3127/NC_O_UNCONNECTED )
  );
  X_BUF   \MASTER/$4I3128/NC  (
    .I(M_CBE4),
    .O(\NLW_MASTER/$4I3128/NC_O_UNCONNECTED )
  );
  X_BUF   \MASTER/$4I3129/NC  (
    .I(M_CBE3),
    .O(\NLW_MASTER/$4I3129/NC_O_UNCONNECTED )
  );
  X_BUF   \MASTER/$4I3130/NC  (
    .I(M_CBE2),
    .O(\NLW_MASTER/$4I3130/NC_O_UNCONNECTED )
  );
  X_BUF   \MASTER/$4I3131/NC  (
    .I(M_CBE1),
    .O(\NLW_MASTER/$4I3131/NC_O_UNCONNECTED )
  );
  X_BUF   \MASTER/$4I3132/NC  (
    .I(M_CBE0),
    .O(\NLW_MASTER/$4I3132/NC_O_UNCONNECTED )
  );
  X_BUF   \MASTER/$4I3134/NC  (
    .I(\ACK64- ),
    .O(\NLW_MASTER/$4I3134/NC_O_UNCONNECTED )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \MASTER/GNT_IOB/IFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(\MASTER/GNT_IOB/$1N2286 ),
    .CLK(CLK),
    .I(GNT_IN),
    .O(\GNT- ),
    .RST(GND)
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \MASTER/GNT_IOB/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(\MASTER/GNT_IOB/$1N2289 ),
    .CLK(CLK),
    .I(\MASTER/NS_GNT- ),
    .O(\MASTER/GNT_O ),
    .RST(GND)
  );
  X_ONE   \MASTER/GNT_IOB/$1I2285/$1I2220  (
    .O(\MASTER/GNT_IOB/$1I2285/$1N2216 )
  );
  X_BUF   \MASTER/GNT_IOB/$1I2285/H  (
    .I(\MASTER/GNT_IOB/$1I2285/$1N2216 ),
    .O(\MASTER/GNT_IOB/$1N2286 )
  );
  X_ONE   \MASTER/GNT_IOB/$1I2288/$1I2220  (
    .O(\MASTER/GNT_IOB/$1I2288/$1N2216 )
  );
  X_BUF   \MASTER/GNT_IOB/$1I2288/H  (
    .I(\MASTER/GNT_IOB/$1I2288/$1N2216 ),
    .O(\MASTER/GNT_IOB/$1N2289 )
  );
  X_ZERO   \MASTER/$4I3148/$1I2218  (
    .O(\MASTER/$4I3148/$1N2216 )
  );
  X_BUF   \MASTER/$4I3148/L  (
    .I(\MASTER/$4I3148/$1N2216 ),
    .O(\MASTER/NS_GNT- )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \MASTER/REQ_IOB/IFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(\MASTER/REQ_IOB/$1N2286 ),
    .CLK(CLK),
    .I(\MASTER/$4N3302 ),
    .O(\MASTER/REQ- ),
    .RST(GND)
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \MASTER/REQ_IOB/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(\MASTER/REQ_IOB/$1N2289 ),
    .CLK(CLK),
    .I(\MASTER/NS_REQ- ),
    .O(REQ_OUT),
    .RST(GND)
  );
  X_ONE   \MASTER/REQ_IOB/$1I2285/$1I2220  (
    .O(\MASTER/REQ_IOB/$1I2285/$1N2216 )
  );
  X_BUF   \MASTER/REQ_IOB/$1I2285/H  (
    .I(\MASTER/REQ_IOB/$1I2285/$1N2216 ),
    .O(\MASTER/REQ_IOB/$1N2286 )
  );
  X_ONE   \MASTER/REQ_IOB/$1I2288/$1I2220  (
    .O(\MASTER/REQ_IOB/$1I2288/$1N2216 )
  );
  X_BUF   \MASTER/REQ_IOB/$1I2288/H  (
    .I(\MASTER/REQ_IOB/$1I2288/$1N2216 ),
    .O(\MASTER/REQ_IOB/$1N2289 )
  );
  X_BUF   \MASTER/$4I3169/NC  (
    .I(\MASTER/REQ- ),
    .O(\NLW_MASTER/$4I3169/NC_O_UNCONNECTED )
  );
  X_AND3   \MASTER/LAT_TIMR/$2I56  (
    .I0(\NlwInverterSignal_MASTER/LAT_TIMR/$2I56/I0 ),
    .I1(\NlwInverterSignal_MASTER/LAT_TIMR/$2I56/I1 ),
    .I2(\NlwInverterSignal_MASTER/LAT_TIMR/$2I56/I2 ),
    .O(\MASTER/LAT_TIMR/T000X )
  );
  X_INV   \MASTER/LAT_TIMR/$2I51  (
    .I(\MASTER/CNT_VAL0 ),
    .O(\MASTER/LAT_TIMR/$2N31 )
  );
  X_AND4   \MASTER/LAT_TIMR/$2I23  (
    .I0(\NlwInverterSignal_MASTER/LAT_TIMR/$2I23/I0 ),
    .I1(\NlwInverterSignal_MASTER/LAT_TIMR/$2I23/I1 ),
    .I2(\NlwInverterSignal_MASTER/LAT_TIMR/$2I23/I2 ),
    .I3(\NlwInverterSignal_MASTER/LAT_TIMR/$2I23/I3 ),
    .O(\MASTER/LAT_TIMR/T4 )
  );
  X_AND3   \MASTER/LAT_TIMR/$2I21  (
    .I0(\NlwInverterSignal_MASTER/LAT_TIMR/$2I21/I0 ),
    .I1(\NlwInverterSignal_MASTER/LAT_TIMR/$2I21/I1 ),
    .I2(\NlwInverterSignal_MASTER/LAT_TIMR/$2I21/I2 ),
    .O(\MASTER/LAT_TIMR/T3 )
  );
  X_AND2   \MASTER/LAT_TIMR/$2I19  (
    .I0(\NlwInverterSignal_MASTER/LAT_TIMR/$2I19/I0 ),
    .I1(\NlwInverterSignal_MASTER/LAT_TIMR/$2I19/I1 ),
    .O(\MASTER/LAT_TIMR/T2 )
  );
  X_AND2   \MASTER/LAT_TIMR/$1I85  (
    .I0(CFG112),
    .I1(\MASTER/LAT_TIMR/TC ),
    .O(\MASTER/LAT_TIMR/$1N74 )
  );
  X_AND3   \MASTER/LAT_TIMR/$1I8  (
    .I0(\NlwInverterSignal_MASTER/LAT_TIMR/$1I8/I0 ),
    .I1(\NlwInverterSignal_MASTER/LAT_TIMR/$1I8/I1 ),
    .I2(\MASTER/LAT_TIMR/T4 ),
    .O(\MASTER/LAT_TIMR/T6 )
  );
  X_INV   \MASTER/LAT_TIMR/$1I71  (
    .I(M_DATA_INT),
    .O(\MASTER/LAT_TIMR/$1N76 )
  );
  X_AND5   \MASTER/LAT_TIMR/$1I29  (
    .I0(\NlwInverterSignal_MASTER/LAT_TIMR/$1I29/I0 ),
    .I1(\NlwInverterSignal_MASTER/LAT_TIMR/$1I29/I1 ),
    .I2(\NlwInverterSignal_MASTER/LAT_TIMR/$1I29/I2 ),
    .I3(\NlwInverterSignal_MASTER/LAT_TIMR/$1I29/I3 ),
    .I4(\MASTER/LAT_TIMR/T000X ),
    .O(\MASTER/LAT_TIMR/TC )
  );
  X_AND4   \MASTER/LAT_TIMR/$1I25  (
    .I0(\NlwInverterSignal_MASTER/LAT_TIMR/$1I25/I0 ),
    .I1(\NlwInverterSignal_MASTER/LAT_TIMR/$1I25/I1 ),
    .I2(\NlwInverterSignal_MASTER/LAT_TIMR/$1I25/I2 ),
    .I3(\MASTER/LAT_TIMR/T4 ),
    .O(\MASTER/LAT_TIMR/T7 )
  );
  X_AND2   \MASTER/LAT_TIMR/$1I11  (
    .I0(\NlwInverterSignal_MASTER/LAT_TIMR/$1I11/I0 ),
    .I1(\MASTER/LAT_TIMR/T4 ),
    .O(\MASTER/LAT_TIMR/T5 )
  );
  X_ONE   \MASTER/LAT_TIMR/$1I129/$1I2220  (
    .O(\MASTER/LAT_TIMR/$1I129/$1N2216 )
  );
  X_BUF   \MASTER/LAT_TIMR/$1I129/H  (
    .I(\MASTER/LAT_TIMR/$1I129/$1N2216 ),
    .O(\MASTER/LAT_TIMR/OR_CE_L )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \MASTER/LAT_TIMR/Q4/$1I35  (
    .CE(\MASTER/LAT_TIMR/OR_CE_L ),
    .CLK(CLK),
    .I(\MASTER/LAT_TIMR/Q4/MD ),
    .O(\MASTER/CNT_VAL4 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \MASTER/LAT_TIMR/Q4/$1I32  (
    .I0(\MASTER/LAT_TIMR/T4 ),
    .I1(\MASTER/CNT_VAL4 ),
    .O(\MASTER/LAT_TIMR/Q4/TQ )
  );
  X_AND2   \MASTER/LAT_TIMR/Q4/$1I30/$1I9  (
    .I0(\MASTER/LAT_TIME4 ),
    .I1(\IFRAME_I- ),
    .O(\MASTER/LAT_TIMR/Q4/$1I30/M1 )
  );
  X_OR2   \MASTER/LAT_TIMR/Q4/$1I30/$1I8  (
    .I0(\MASTER/LAT_TIMR/Q4/$1I30/M1 ),
    .I1(\MASTER/LAT_TIMR/Q4/$1I30/M0 ),
    .O(\MASTER/LAT_TIMR/Q4/MD )
  );
  X_AND2   \MASTER/LAT_TIMR/Q4/$1I30/$1I7  (
    .I0(\NlwInverterSignal_MASTER/LAT_TIMR/Q4/$1I30/$1I7/I0 ),
    .I1(\MASTER/LAT_TIMR/Q4/TQ ),
    .O(\MASTER/LAT_TIMR/Q4/$1I30/M0 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \MASTER/LAT_TIMR/Q6/$1I35  (
    .CE(\MASTER/LAT_TIMR/OR_CE_L ),
    .CLK(CLK),
    .I(\MASTER/LAT_TIMR/Q6/MD ),
    .O(\MASTER/CNT_VAL6 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \MASTER/LAT_TIMR/Q6/$1I32  (
    .I0(\MASTER/LAT_TIMR/T6 ),
    .I1(\MASTER/CNT_VAL6 ),
    .O(\MASTER/LAT_TIMR/Q6/TQ )
  );
  X_AND2   \MASTER/LAT_TIMR/Q6/$1I30/$1I9  (
    .I0(\MASTER/LAT_TIME6 ),
    .I1(\IFRAME_I- ),
    .O(\MASTER/LAT_TIMR/Q6/$1I30/M1 )
  );
  X_OR2   \MASTER/LAT_TIMR/Q6/$1I30/$1I8  (
    .I0(\MASTER/LAT_TIMR/Q6/$1I30/M1 ),
    .I1(\MASTER/LAT_TIMR/Q6/$1I30/M0 ),
    .O(\MASTER/LAT_TIMR/Q6/MD )
  );
  X_AND2   \MASTER/LAT_TIMR/Q6/$1I30/$1I7  (
    .I0(\NlwInverterSignal_MASTER/LAT_TIMR/Q6/$1I30/$1I7/I0 ),
    .I1(\MASTER/LAT_TIMR/Q6/TQ ),
    .O(\MASTER/LAT_TIMR/Q6/$1I30/M0 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \MASTER/LAT_TIMR/Q7/$1I35  (
    .CE(\MASTER/LAT_TIMR/OR_CE_L ),
    .CLK(CLK),
    .I(\MASTER/LAT_TIMR/Q7/MD ),
    .O(\MASTER/CNT_VAL7 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \MASTER/LAT_TIMR/Q7/$1I32  (
    .I0(\MASTER/LAT_TIMR/T7 ),
    .I1(\MASTER/CNT_VAL7 ),
    .O(\MASTER/LAT_TIMR/Q7/TQ )
  );
  X_AND2   \MASTER/LAT_TIMR/Q7/$1I30/$1I9  (
    .I0(\MASTER/LAT_TIME7 ),
    .I1(\IFRAME_I- ),
    .O(\MASTER/LAT_TIMR/Q7/$1I30/M1 )
  );
  X_OR2   \MASTER/LAT_TIMR/Q7/$1I30/$1I8  (
    .I0(\MASTER/LAT_TIMR/Q7/$1I30/M1 ),
    .I1(\MASTER/LAT_TIMR/Q7/$1I30/M0 ),
    .O(\MASTER/LAT_TIMR/Q7/MD )
  );
  X_AND2   \MASTER/LAT_TIMR/Q7/$1I30/$1I7  (
    .I0(\NlwInverterSignal_MASTER/LAT_TIMR/Q7/$1I30/$1I7/I0 ),
    .I1(\MASTER/LAT_TIMR/Q7/TQ ),
    .O(\MASTER/LAT_TIMR/Q7/$1I30/M0 )
  );
  X_AND2   \MASTER/LAT_TIMR/TIME_OUT/$1I2214  (
    .I0(\NlwInverterSignal_MASTER/LAT_TIMR/TIME_OUT/$1I2214/I0 ),
    .I1(NlwRenamedSig_OI_TIME_OUT),
    .O(\MASTER/LAT_TIMR/TIME_OUT/$1N2215 )
  );
  X_OR2   \MASTER/LAT_TIMR/TIME_OUT/$1I2213  (
    .I0(\MASTER/LAT_TIMR/$1N74 ),
    .I1(\MASTER/LAT_TIMR/TIME_OUT/$1N2215 ),
    .O(\MASTER/LAT_TIMR/TIME_OUT/D )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \MASTER/LAT_TIMR/TIME_OUT/FDCE  (
    .CE(VCC),
    .CLK(CLK),
    .I(\MASTER/LAT_TIMR/TIME_OUT/D ),
    .O(NlwRenamedSig_OI_TIME_OUT),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \MASTER/LAT_TIMR/Q5/$1I35  (
    .CE(\MASTER/LAT_TIMR/OR_CE_L ),
    .CLK(CLK),
    .I(\MASTER/LAT_TIMR/Q5/MD ),
    .O(\MASTER/CNT_VAL5 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \MASTER/LAT_TIMR/Q5/$1I32  (
    .I0(\MASTER/LAT_TIMR/T5 ),
    .I1(\MASTER/CNT_VAL5 ),
    .O(\MASTER/LAT_TIMR/Q5/TQ )
  );
  X_AND2   \MASTER/LAT_TIMR/Q5/$1I30/$1I9  (
    .I0(\MASTER/LAT_TIME5 ),
    .I1(\IFRAME_I- ),
    .O(\MASTER/LAT_TIMR/Q5/$1I30/M1 )
  );
  X_OR2   \MASTER/LAT_TIMR/Q5/$1I30/$1I8  (
    .I0(\MASTER/LAT_TIMR/Q5/$1I30/M1 ),
    .I1(\MASTER/LAT_TIMR/Q5/$1I30/M0 ),
    .O(\MASTER/LAT_TIMR/Q5/MD )
  );
  X_AND2   \MASTER/LAT_TIMR/Q5/$1I30/$1I7  (
    .I0(\NlwInverterSignal_MASTER/LAT_TIMR/Q5/$1I30/$1I7/I0 ),
    .I1(\MASTER/LAT_TIMR/Q5/TQ ),
    .O(\MASTER/LAT_TIMR/Q5/$1I30/M0 )
  );
  X_ONE   \MASTER/LAT_TIMR/$2I121/$1I2220  (
    .O(\MASTER/LAT_TIMR/$2I121/$1N2216 )
  );
  X_BUF   \MASTER/LAT_TIMR/$2I121/H  (
    .I(\MASTER/LAT_TIMR/$2I121/$1N2216 ),
    .O(\MASTER/LAT_TIMR/$2N13 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \MASTER/LAT_TIMR/Q1/$1I35  (
    .CE(\MASTER/LAT_TIMR/OR_CE_L ),
    .CLK(CLK),
    .I(\MASTER/LAT_TIMR/Q1/MD ),
    .O(\MASTER/CNT_VAL1 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \MASTER/LAT_TIMR/Q1/$1I32  (
    .I0(\MASTER/LAT_TIMR/$2N31 ),
    .I1(\MASTER/CNT_VAL1 ),
    .O(\MASTER/LAT_TIMR/Q1/TQ )
  );
  X_AND2   \MASTER/LAT_TIMR/Q1/$1I30/$1I9  (
    .I0(\MASTER/LAT_TIME1 ),
    .I1(\IFRAME_I- ),
    .O(\MASTER/LAT_TIMR/Q1/$1I30/M1 )
  );
  X_OR2   \MASTER/LAT_TIMR/Q1/$1I30/$1I8  (
    .I0(\MASTER/LAT_TIMR/Q1/$1I30/M1 ),
    .I1(\MASTER/LAT_TIMR/Q1/$1I30/M0 ),
    .O(\MASTER/LAT_TIMR/Q1/MD )
  );
  X_AND2   \MASTER/LAT_TIMR/Q1/$1I30/$1I7  (
    .I0(\NlwInverterSignal_MASTER/LAT_TIMR/Q1/$1I30/$1I7/I0 ),
    .I1(\MASTER/LAT_TIMR/Q1/TQ ),
    .O(\MASTER/LAT_TIMR/Q1/$1I30/M0 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \MASTER/LAT_TIMR/Q0/$1I35  (
    .CE(\MASTER/LAT_TIMR/OR_CE_L ),
    .CLK(CLK),
    .I(\MASTER/LAT_TIMR/Q0/MD ),
    .O(\MASTER/CNT_VAL0 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \MASTER/LAT_TIMR/Q0/$1I32  (
    .I0(\MASTER/LAT_TIMR/$2N13 ),
    .I1(\MASTER/CNT_VAL0 ),
    .O(\MASTER/LAT_TIMR/Q0/TQ )
  );
  X_AND2   \MASTER/LAT_TIMR/Q0/$1I30/$1I9  (
    .I0(\MASTER/LAT_TIME0 ),
    .I1(\IFRAME_I- ),
    .O(\MASTER/LAT_TIMR/Q0/$1I30/M1 )
  );
  X_OR2   \MASTER/LAT_TIMR/Q0/$1I30/$1I8  (
    .I0(\MASTER/LAT_TIMR/Q0/$1I30/M1 ),
    .I1(\MASTER/LAT_TIMR/Q0/$1I30/M0 ),
    .O(\MASTER/LAT_TIMR/Q0/MD )
  );
  X_AND2   \MASTER/LAT_TIMR/Q0/$1I30/$1I7  (
    .I0(\NlwInverterSignal_MASTER/LAT_TIMR/Q0/$1I30/$1I7/I0 ),
    .I1(\MASTER/LAT_TIMR/Q0/TQ ),
    .O(\MASTER/LAT_TIMR/Q0/$1I30/M0 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \MASTER/LAT_TIMR/Q2/$1I35  (
    .CE(\MASTER/LAT_TIMR/OR_CE_L ),
    .CLK(CLK),
    .I(\MASTER/LAT_TIMR/Q2/MD ),
    .O(\MASTER/CNT_VAL2 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \MASTER/LAT_TIMR/Q2/$1I32  (
    .I0(\MASTER/LAT_TIMR/T2 ),
    .I1(\MASTER/CNT_VAL2 ),
    .O(\MASTER/LAT_TIMR/Q2/TQ )
  );
  X_AND2   \MASTER/LAT_TIMR/Q2/$1I30/$1I9  (
    .I0(\MASTER/LAT_TIME2 ),
    .I1(\IFRAME_I- ),
    .O(\MASTER/LAT_TIMR/Q2/$1I30/M1 )
  );
  X_OR2   \MASTER/LAT_TIMR/Q2/$1I30/$1I8  (
    .I0(\MASTER/LAT_TIMR/Q2/$1I30/M1 ),
    .I1(\MASTER/LAT_TIMR/Q2/$1I30/M0 ),
    .O(\MASTER/LAT_TIMR/Q2/MD )
  );
  X_AND2   \MASTER/LAT_TIMR/Q2/$1I30/$1I7  (
    .I0(\NlwInverterSignal_MASTER/LAT_TIMR/Q2/$1I30/$1I7/I0 ),
    .I1(\MASTER/LAT_TIMR/Q2/TQ ),
    .O(\MASTER/LAT_TIMR/Q2/$1I30/M0 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \MASTER/LAT_TIMR/Q3/$1I35  (
    .CE(\MASTER/LAT_TIMR/OR_CE_L ),
    .CLK(CLK),
    .I(\MASTER/LAT_TIMR/Q3/MD ),
    .O(\MASTER/CNT_VAL3 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \MASTER/LAT_TIMR/Q3/$1I32  (
    .I0(\MASTER/LAT_TIMR/T3 ),
    .I1(\MASTER/CNT_VAL3 ),
    .O(\MASTER/LAT_TIMR/Q3/TQ )
  );
  X_AND2   \MASTER/LAT_TIMR/Q3/$1I30/$1I9  (
    .I0(\MASTER/LAT_TIME3 ),
    .I1(\IFRAME_I- ),
    .O(\MASTER/LAT_TIMR/Q3/$1I30/M1 )
  );
  X_OR2   \MASTER/LAT_TIMR/Q3/$1I30/$1I8  (
    .I0(\MASTER/LAT_TIMR/Q3/$1I30/M1 ),
    .I1(\MASTER/LAT_TIMR/Q3/$1I30/M0 ),
    .O(\MASTER/LAT_TIMR/Q3/MD )
  );
  X_AND2   \MASTER/LAT_TIMR/Q3/$1I30/$1I7  (
    .I0(\NlwInverterSignal_MASTER/LAT_TIMR/Q3/$1I30/$1I7/I0 ),
    .I1(\MASTER/LAT_TIMR/Q3/TQ ),
    .O(\MASTER/LAT_TIMR/Q3/$1I30/M0 )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2526  (
    .I(\MASTER/PCI-0CH/$1N2518 ),
    .O(\MASTER/REG_0CH0 )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2525  (
    .I(\MASTER/PCI-0CH/$1N2518 ),
    .O(\MASTER/REG_0CH1 )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2524  (
    .I(\MASTER/PCI-0CH/$1N2518 ),
    .O(\MASTER/REG_0CH2 )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2523  (
    .I(\MASTER/PCI-0CH/$1N2518 ),
    .O(\MASTER/REG_0CH3 )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2522  (
    .I(\MASTER/PCI-0CH/$1N2518 ),
    .O(\MASTER/REG_0CH4 )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2521  (
    .I(\MASTER/PCI-0CH/$1N2518 ),
    .O(\MASTER/REG_0CH5 )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2520  (
    .I(\MASTER/PCI-0CH/$1N2518 ),
    .O(\MASTER/REG_0CH6 )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2519  (
    .I(\MASTER/PCI-0CH/$1N2518 ),
    .O(\MASTER/REG_0CH7 )
  );
  X_ZERO   \MASTER/PCI-0CH/$1I2517  (
    .O(\MASTER/PCI-0CH/$1N2518 )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2512  (
    .I(\MASTER/PCI-0CH/$1N2513 ),
    .O(\MASTER/REG_0CH16 )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2511  (
    .I(\MASTER/PCI-0CH/$1N2513 ),
    .O(\MASTER/REG_0CH17 )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2510  (
    .I(\MASTER/PCI-0CH/$1N2513 ),
    .O(\MASTER/REG_0CH18 )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2509  (
    .I(\MASTER/PCI-0CH/$1N2513 ),
    .O(\MASTER/REG_0CH19 )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2508  (
    .I(\MASTER/PCI-0CH/$1N2513 ),
    .O(\MASTER/REG_0CH20 )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2507  (
    .I(\MASTER/PCI-0CH/$1N2513 ),
    .O(\MASTER/REG_0CH21 )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2506  (
    .I(\MASTER/PCI-0CH/$1N2513 ),
    .O(\MASTER/REG_0CH22 )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2505  (
    .I(\MASTER/PCI-0CH/$1N2513 ),
    .O(\MASTER/REG_0CH23 )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2504  (
    .I(\MASTER/PCI-0CH/$1N2513 ),
    .O(\MASTER/REG_0CH24 )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2503  (
    .I(\MASTER/PCI-0CH/$1N2513 ),
    .O(\MASTER/REG_0CH25 )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2502  (
    .I(\MASTER/PCI-0CH/$1N2513 ),
    .O(\MASTER/REG_0CH26 )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2501  (
    .I(\MASTER/PCI-0CH/$1N2513 ),
    .O(\MASTER/REG_0CH27 )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2500  (
    .I(\MASTER/PCI-0CH/$1N2513 ),
    .O(\MASTER/REG_0CH28 )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2499  (
    .I(\MASTER/PCI-0CH/$1N2513 ),
    .O(\MASTER/REG_0CH29 )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2498  (
    .I(\MASTER/PCI-0CH/$1N2513 ),
    .O(\MASTER/REG_0CH30 )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2497  (
    .I(\MASTER/PCI-0CH/$1N2513 ),
    .O(\MASTER/REG_0CH31 )
  );
  X_ZERO   \MASTER/PCI-0CH/$1I2493  (
    .O(\MASTER/PCI-0CH/$1N2513 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \MASTER/PCI-0CH/LAT-TIME/Q7  (
    .CE(CE3_1),
    .CLK(CLK),
    .I(ADIO15),
    .O(\MASTER/REG_0CH15 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \MASTER/PCI-0CH/LAT-TIME/Q1  (
    .CE(CE3_1),
    .CLK(CLK),
    .I(ADIO9),
    .O(\MASTER/REG_0CH9 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \MASTER/PCI-0CH/LAT-TIME/Q5  (
    .CE(CE3_1),
    .CLK(CLK),
    .I(ADIO13),
    .O(\MASTER/REG_0CH13 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \MASTER/PCI-0CH/LAT-TIME/Q3  (
    .CE(CE3_1),
    .CLK(CLK),
    .I(ADIO11),
    .O(\MASTER/REG_0CH11 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \MASTER/PCI-0CH/LAT-TIME/Q0  (
    .CE(CE3_1),
    .CLK(CLK),
    .I(ADIO8),
    .O(\MASTER/REG_0CH8 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \MASTER/PCI-0CH/LAT-TIME/Q2  (
    .CE(CE3_1),
    .CLK(CLK),
    .I(ADIO10),
    .O(\MASTER/REG_0CH10 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \MASTER/PCI-0CH/LAT-TIME/Q4  (
    .CE(CE3_1),
    .CLK(CLK),
    .I(ADIO12),
    .O(\MASTER/REG_0CH12 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \MASTER/PCI-0CH/LAT-TIME/Q6  (
    .CE(CE3_1),
    .CLK(CLK),
    .I(ADIO14),
    .O(\MASTER/REG_0CH14 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_BUF   \MASTER/PCI-0CH/$1I2529/NC  (
    .I(CE3_2),
    .O(\NLW_MASTER/PCI-0CH/$1I2529/NC_O_UNCONNECTED )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2532/NC  (
    .I(CE3_0),
    .O(\NLW_MASTER/PCI-0CH/$1I2532/NC_O_UNCONNECTED )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2534/NC  (
    .I(CE3_3),
    .O(\NLW_MASTER/PCI-0CH/$1I2534/NC_O_UNCONNECTED )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2536/NC  (
    .I(ADIO31),
    .O(\NLW_MASTER/PCI-0CH/$1I2536/NC_O_UNCONNECTED )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2538/NC  (
    .I(ADIO30),
    .O(\NLW_MASTER/PCI-0CH/$1I2538/NC_O_UNCONNECTED )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2540/NC  (
    .I(ADIO29),
    .O(\NLW_MASTER/PCI-0CH/$1I2540/NC_O_UNCONNECTED )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2542/NC  (
    .I(ADIO28),
    .O(\NLW_MASTER/PCI-0CH/$1I2542/NC_O_UNCONNECTED )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2544/NC  (
    .I(ADIO27),
    .O(\NLW_MASTER/PCI-0CH/$1I2544/NC_O_UNCONNECTED )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2546/NC  (
    .I(ADIO26),
    .O(\NLW_MASTER/PCI-0CH/$1I2546/NC_O_UNCONNECTED )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2548/NC  (
    .I(ADIO25),
    .O(\NLW_MASTER/PCI-0CH/$1I2548/NC_O_UNCONNECTED )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2550/NC  (
    .I(ADIO24),
    .O(\NLW_MASTER/PCI-0CH/$1I2550/NC_O_UNCONNECTED )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2552/NC  (
    .I(ADIO23),
    .O(\NLW_MASTER/PCI-0CH/$1I2552/NC_O_UNCONNECTED )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2554/NC  (
    .I(ADIO22),
    .O(\NLW_MASTER/PCI-0CH/$1I2554/NC_O_UNCONNECTED )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2556/NC  (
    .I(ADIO21),
    .O(\NLW_MASTER/PCI-0CH/$1I2556/NC_O_UNCONNECTED )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2558/NC  (
    .I(ADIO20),
    .O(\NLW_MASTER/PCI-0CH/$1I2558/NC_O_UNCONNECTED )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2560/NC  (
    .I(ADIO19),
    .O(\NLW_MASTER/PCI-0CH/$1I2560/NC_O_UNCONNECTED )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2562/NC  (
    .I(ADIO18),
    .O(\NLW_MASTER/PCI-0CH/$1I2562/NC_O_UNCONNECTED )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2564/NC  (
    .I(ADIO17),
    .O(\NLW_MASTER/PCI-0CH/$1I2564/NC_O_UNCONNECTED )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2566/NC  (
    .I(ADIO16),
    .O(\NLW_MASTER/PCI-0CH/$1I2566/NC_O_UNCONNECTED )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2568/NC  (
    .I(ADIO7),
    .O(\NLW_MASTER/PCI-0CH/$1I2568/NC_O_UNCONNECTED )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2570/NC  (
    .I(ADIO6),
    .O(\NLW_MASTER/PCI-0CH/$1I2570/NC_O_UNCONNECTED )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2572/NC  (
    .I(ADIO5),
    .O(\NLW_MASTER/PCI-0CH/$1I2572/NC_O_UNCONNECTED )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2574/NC  (
    .I(ADIO4),
    .O(\NLW_MASTER/PCI-0CH/$1I2574/NC_O_UNCONNECTED )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2576/NC  (
    .I(ADIO3),
    .O(\NLW_MASTER/PCI-0CH/$1I2576/NC_O_UNCONNECTED )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2578/NC  (
    .I(ADIO2),
    .O(\NLW_MASTER/PCI-0CH/$1I2578/NC_O_UNCONNECTED )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2580/NC  (
    .I(ADIO1),
    .O(\NLW_MASTER/PCI-0CH/$1I2580/NC_O_UNCONNECTED )
  );
  X_BUF   \MASTER/PCI-0CH/$1I2582/NC  (
    .I(ADIO0),
    .O(\NLW_MASTER/PCI-0CH/$1I2582/NC_O_UNCONNECTED )
  );
  X_TRI   \MASTER/3/UPPER/T0  (
    .I(\MASTER/REG_0CH16 ),
    .O(ADIO16),
    .CTL(\NlwInverterSignal_MASTER/3/UPPER/T0/T )
  );
  X_TRI   \MASTER/3/UPPER/T1  (
    .I(\MASTER/REG_0CH17 ),
    .O(ADIO17),
    .CTL(\NlwInverterSignal_MASTER/3/UPPER/T1/T )
  );
  X_TRI   \MASTER/3/UPPER/T2  (
    .I(\MASTER/REG_0CH18 ),
    .O(ADIO18),
    .CTL(\NlwInverterSignal_MASTER/3/UPPER/T2/T )
  );
  X_TRI   \MASTER/3/UPPER/T3  (
    .I(\MASTER/REG_0CH19 ),
    .O(ADIO19),
    .CTL(\NlwInverterSignal_MASTER/3/UPPER/T3/T )
  );
  X_TRI   \MASTER/3/UPPER/T4  (
    .I(\MASTER/REG_0CH20 ),
    .O(ADIO20),
    .CTL(\NlwInverterSignal_MASTER/3/UPPER/T4/T )
  );
  X_TRI   \MASTER/3/UPPER/T5  (
    .I(\MASTER/REG_0CH21 ),
    .O(ADIO21),
    .CTL(\NlwInverterSignal_MASTER/3/UPPER/T5/T )
  );
  X_TRI   \MASTER/3/UPPER/T6  (
    .I(\MASTER/REG_0CH22 ),
    .O(ADIO22),
    .CTL(\NlwInverterSignal_MASTER/3/UPPER/T6/T )
  );
  X_TRI   \MASTER/3/UPPER/T7  (
    .I(\MASTER/REG_0CH23 ),
    .O(ADIO23),
    .CTL(\NlwInverterSignal_MASTER/3/UPPER/T7/T )
  );
  X_TRI   \MASTER/3/UPPER/T8  (
    .I(\MASTER/REG_0CH24 ),
    .O(ADIO24),
    .CTL(\NlwInverterSignal_MASTER/3/UPPER/T8/T )
  );
  X_TRI   \MASTER/3/UPPER/T9  (
    .I(\MASTER/REG_0CH25 ),
    .O(ADIO25),
    .CTL(\NlwInverterSignal_MASTER/3/UPPER/T9/T )
  );
  X_TRI   \MASTER/3/UPPER/T10  (
    .I(\MASTER/REG_0CH26 ),
    .O(ADIO26),
    .CTL(\NlwInverterSignal_MASTER/3/UPPER/T10/T )
  );
  X_TRI   \MASTER/3/UPPER/T11  (
    .I(\MASTER/REG_0CH27 ),
    .O(ADIO27),
    .CTL(\NlwInverterSignal_MASTER/3/UPPER/T11/T )
  );
  X_TRI   \MASTER/3/UPPER/T12  (
    .I(\MASTER/REG_0CH28 ),
    .O(ADIO28),
    .CTL(\NlwInverterSignal_MASTER/3/UPPER/T12/T )
  );
  X_TRI   \MASTER/3/UPPER/T13  (
    .I(\MASTER/REG_0CH29 ),
    .O(ADIO29),
    .CTL(\NlwInverterSignal_MASTER/3/UPPER/T13/T )
  );
  X_TRI   \MASTER/3/UPPER/T14  (
    .I(\MASTER/REG_0CH30 ),
    .O(ADIO30),
    .CTL(\NlwInverterSignal_MASTER/3/UPPER/T14/T )
  );
  X_TRI   \MASTER/3/UPPER/T15  (
    .I(\MASTER/REG_0CH31 ),
    .O(ADIO31),
    .CTL(\NlwInverterSignal_MASTER/3/UPPER/T15/T )
  );
  X_TRI   \MASTER/3/LOWER/T0  (
    .I(\MASTER/REG_0CH0 ),
    .O(ADIO0),
    .CTL(\NlwInverterSignal_MASTER/3/LOWER/T0/T )
  );
  X_TRI   \MASTER/3/LOWER/T1  (
    .I(\MASTER/REG_0CH1 ),
    .O(ADIO1),
    .CTL(\NlwInverterSignal_MASTER/3/LOWER/T1/T )
  );
  X_TRI   \MASTER/3/LOWER/T2  (
    .I(\MASTER/REG_0CH2 ),
    .O(ADIO2),
    .CTL(\NlwInverterSignal_MASTER/3/LOWER/T2/T )
  );
  X_TRI   \MASTER/3/LOWER/T3  (
    .I(\MASTER/REG_0CH3 ),
    .O(ADIO3),
    .CTL(\NlwInverterSignal_MASTER/3/LOWER/T3/T )
  );
  X_TRI   \MASTER/3/LOWER/T4  (
    .I(\MASTER/REG_0CH4 ),
    .O(ADIO4),
    .CTL(\NlwInverterSignal_MASTER/3/LOWER/T4/T )
  );
  X_TRI   \MASTER/3/LOWER/T5  (
    .I(\MASTER/REG_0CH5 ),
    .O(ADIO5),
    .CTL(\NlwInverterSignal_MASTER/3/LOWER/T5/T )
  );
  X_TRI   \MASTER/3/LOWER/T6  (
    .I(\MASTER/REG_0CH6 ),
    .O(ADIO6),
    .CTL(\NlwInverterSignal_MASTER/3/LOWER/T6/T )
  );
  X_TRI   \MASTER/3/LOWER/T7  (
    .I(\MASTER/REG_0CH7 ),
    .O(ADIO7),
    .CTL(\NlwInverterSignal_MASTER/3/LOWER/T7/T )
  );
  X_TRI   \MASTER/3/LOWER/T8  (
    .I(\MASTER/REG_0CH8 ),
    .O(ADIO8),
    .CTL(\NlwInverterSignal_MASTER/3/LOWER/T8/T )
  );
  X_TRI   \MASTER/3/LOWER/T9  (
    .I(\MASTER/REG_0CH9 ),
    .O(ADIO9),
    .CTL(\NlwInverterSignal_MASTER/3/LOWER/T9/T )
  );
  X_TRI   \MASTER/3/LOWER/T10  (
    .I(\MASTER/REG_0CH10 ),
    .O(ADIO10),
    .CTL(\NlwInverterSignal_MASTER/3/LOWER/T10/T )
  );
  X_TRI   \MASTER/3/LOWER/T11  (
    .I(\MASTER/REG_0CH11 ),
    .O(ADIO11),
    .CTL(\NlwInverterSignal_MASTER/3/LOWER/T11/T )
  );
  X_TRI   \MASTER/3/LOWER/T12  (
    .I(\MASTER/REG_0CH12 ),
    .O(ADIO12),
    .CTL(\NlwInverterSignal_MASTER/3/LOWER/T12/T )
  );
  X_TRI   \MASTER/3/LOWER/T13  (
    .I(\MASTER/REG_0CH13 ),
    .O(ADIO13),
    .CTL(\NlwInverterSignal_MASTER/3/LOWER/T13/T )
  );
  X_TRI   \MASTER/3/LOWER/T14  (
    .I(\MASTER/REG_0CH14 ),
    .O(ADIO14),
    .CTL(\NlwInverterSignal_MASTER/3/LOWER/T14/T )
  );
  X_TRI   \MASTER/3/LOWER/T15  (
    .I(\MASTER/REG_0CH15 ),
    .O(ADIO15),
    .CTL(\NlwInverterSignal_MASTER/3/LOWER/T15/T )
  );
  X_BUF   \MASTER/$4I3247/NC  (
    .I(\MASTER/IREQ- ),
    .O(\NLW_MASTER/$4I3247/NC_O_UNCONNECTED )
  );
  X_ZERO   \MASTER/$4I3254/$1I2218  (
    .O(\MASTER/$4I3254/$1N2216 )
  );
  X_BUF   \MASTER/$4I3254/L  (
    .I(\MASTER/$4I3254/$1N2216 ),
    .O(\MASTER/$4N3252 )
  );
  X_BUF   \MASTER/$4I3298/NC  (
    .I(\MASTER/IREQ64- ),
    .O(\NLW_MASTER/$4I3298/NC_O_UNCONNECTED )
  );
  X_BUF   \MASTER/$4I3318/NC  (
    .I(\MASTER/GNT_O ),
    .O(\NLW_MASTER/$4I3318/NC_O_UNCONNECTED )
  );
  X_ONE   \MASTER/$4I3319/$1I2220  (
    .O(\MASTER/$4I3319/$1N2216 )
  );
  X_BUF   \MASTER/$4I3319/H  (
    .I(\MASTER/$4I3319/$1N2216 ),
    .O(\MASTER/$4N3302 )
  );
  X_OR2   \PCI-CNTL/$4I804  (
    .I0(BACKOFF_INT),
    .I1(S_DATA_INT),
    .O(\PCI-CNTL/HOLDCYC )
  );
  X_AND3   \PCI-CNTL/$4I788  (
    .I0(\NlwInverterSignal_PCI-CNTL/$4I788/I0 ),
    .I1(S_DATA_INT),
    .I2(NlwRenamedSig_OI_S_WRDN),
    .O(\PCI-CNTL/WIN_3628 )
  );
  X_OR2   \PCI-CNTL/$4I749  (
    .I0(\PCI-CNTL/ANY_BH64 ),
    .I1(\PCI-CNTL/ANY_NS_BH64 ),
    .O(\PCI-CNTL/$4N752 )
  );
  X_OR3   \PCI-CNTL/$4I738  (
    .I0(BH64_2),
    .I1(BH64_1),
    .I2(BH64_0),
    .O(\PCI-CNTL/ANY_BH64 )
  );
  X_OR3   \PCI-CNTL/$4I736  (
    .I0(NS_BH64_2),
    .I1(NS_BH64_1),
    .I2(NS_BH64_0),
    .O(\PCI-CNTL/ANY_NS_BH64 )
  );
  X_AND3   \PCI-CNTL/$4I719  (
    .I0(\NlwInverterSignal_PCI-CNTL/$4I719/I0 ),
    .I1(\PCI-CNTL/WIN_3628 ),
    .I2(S_CYCLE64_INT),
    .O(\PCI-CNTL/NS_PWIN64 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PWIN64_FF  (
    .CE(VCC),
    .CLK(CLK),
    .I(\PCI-CNTL/NS_PWIN64 ),
    .O(TPWIN64),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/CYC64_FF  (
    .CE(VCC),
    .CLK(CLK),
    .I(\PCI-CNTL/NS_CYC64 ),
    .O(S_CYCLE64_INT),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PWIN_FF  (
    .CE(VCC),
    .CLK(CLK),
    .I(\PCI-CNTL/NS_PWIN ),
    .O(TPWIN),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND2   \PCI-CNTL/$4I446  (
    .I0(\NlwInverterSignal_PCI-CNTL/$4I446/I0 ),
    .I1(\PCI-CNTL/WIN_3628 ),
    .O(\PCI-CNTL/NS_PWIN )
  );
  X_INV   \PCI-CNTL/$1I999  (
    .I(APERR_N),
    .O(\PCI-CNTL/$1N1000 )
  );
  X_OR2   \PCI-CNTL/$1I985  (
    .I0(BACKOFF_INT),
    .I1(S_DATA_INT),
    .O(\PCI-CNTL/$1N988 )
  );
  X_AND2   \PCI-CNTL/$1I978  (
    .I0(\PCI-CNTL/S_ABORT ),
    .I1(\PCI-CNTL/$1N988 ),
    .O(SET11)
  );
  X_INV   \PCI-CNTL/$1I915  (
    .I(CBE_IN0),
    .O(\PCI-CNTL/CBE_N0 )
  );
  X_INV   \PCI-CNTL/$1I914  (
    .I(CBE_IN1),
    .O(\PCI-CNTL/CBE_N1 )
  );
  X_INV   \PCI-CNTL/$1I913  (
    .I(CBE_IN2),
    .O(\PCI-CNTL/CBE_N2 )
  );
  X_INV   \PCI-CNTL/$1I912  (
    .I(CBE_IN3),
    .O(\PCI-CNTL/CBE_N3 )
  );
  X_AND3   \PCI-CNTL/$1I840  (
    .I0(\NlwInverterSignal_PCI-CNTL/$1I840/I0 ),
    .I1(\NlwInverterSignal_PCI-CNTL/$1I840/I1 ),
    .I2(NlwRenamedSig_OI_S_WRDN),
    .O(\PCI-CNTL/DSTR )
  );
  X_AND2   \PCI-CNTL/$1I823  (
    .I0(\NlwInverterSignal_PCI-CNTL/$1I823/I0 ),
    .I1(\TDEVSEL_I- ),
    .O(\PCI-CNTL/END )
  );
  X_OR3   \PCI-CNTL/$1I1005  (
    .I0(\NlwInverterSignal_PCI-CNTL/$1I1005/I0 ),
    .I1(\PCI-CNTL/HOLD_APERR ),
    .I2(S_ABORT),
    .O(\PCI-CNTL/S_ABORT )
  );
  X_AND2   \PCI-CNTL/PCI-LA/$1I2751  (
    .I0(\PCI-CNTL/PCI-LA/AD7610-0000 ),
    .I1(\PCI-CNTL/PCI-LA/$1N2666 ),
    .O(\PCI-CNTL/ADX0 )
  );
  X_AND2   \PCI-CNTL/PCI-LA/$1I2748  (
    .I0(\PCI-CNTL/PCI-LA/AD7610-0000 ),
    .I1(\PCI-CNTL/PCI-LA/$1N2762 ),
    .O(\PCI-CNTL/ADX1 )
  );
  X_AND2   \PCI-CNTL/PCI-LA/$1I2745  (
    .I0(\PCI-CNTL/PCI-LA/AD7610-0000 ),
    .I1(\PCI-CNTL/PCI-LA/$1N2668 ),
    .O(\PCI-CNTL/ADX2 )
  );
  X_AND2   \PCI-CNTL/PCI-LA/$1I2742  (
    .I0(\PCI-CNTL/PCI-LA/AD7610-0000 ),
    .I1(\PCI-CNTL/PCI-LA/$1N2764 ),
    .O(\PCI-CNTL/ADX3 )
  );
  X_AND2   \PCI-CNTL/PCI-LA/$1I2739  (
    .I0(\PCI-CNTL/PCI-LA/AD7610-0000 ),
    .I1(\PCI-CNTL/PCI-LA/$1N2670 ),
    .O(\PCI-CNTL/ADX4 )
  );
  X_AND2   \PCI-CNTL/PCI-LA/$1I2736  (
    .I0(\PCI-CNTL/PCI-LA/AD7610-0000 ),
    .I1(\PCI-CNTL/PCI-LA/$1N2766 ),
    .O(\PCI-CNTL/ADX5 )
  );
  X_AND2   \PCI-CNTL/PCI-LA/$1I2733  (
    .I0(\PCI-CNTL/PCI-LA/AD7610-0000 ),
    .I1(\PCI-CNTL/PCI-LA/$1N2672 ),
    .O(\PCI-CNTL/ADX6 )
  );
  X_AND2   \PCI-CNTL/PCI-LA/$1I2730  (
    .I0(\PCI-CNTL/PCI-LA/AD7610-0000 ),
    .I1(\PCI-CNTL/PCI-LA/$1N2768 ),
    .O(\PCI-CNTL/ADX7 )
  );
  X_AND2   \PCI-CNTL/PCI-LA/$1I2723  (
    .I0(\PCI-CNTL/PCI-LA/AD7610-0000 ),
    .I1(\PCI-CNTL/PCI-LA/$1N2760 ),
    .O(\PCI-CNTL/ADX8 )
  );
  X_AND2   \PCI-CNTL/PCI-LA/$1I2720  (
    .I0(\PCI-CNTL/PCI-LA/AD7610-0000 ),
    .I1(\PCI-CNTL/PCI-LA/$1N2625 ),
    .O(\PCI-CNTL/ADX9 )
  );
  X_AND2   \PCI-CNTL/PCI-LA/$1I2717  (
    .I0(\PCI-CNTL/PCI-LA/AD7610-0000 ),
    .I1(\PCI-CNTL/PCI-LA/$1N2624 ),
    .O(\PCI-CNTL/ADX10 )
  );
  X_AND2   \PCI-CNTL/PCI-LA/$1I2714  (
    .I0(\PCI-CNTL/PCI-LA/AD7610-0000 ),
    .I1(\PCI-CNTL/PCI-LA/$1N2623 ),
    .O(\PCI-CNTL/ADX11 )
  );
  X_AND2   \PCI-CNTL/PCI-LA/$1I2711  (
    .I0(\PCI-CNTL/PCI-LA/AD7610-0000 ),
    .I1(\PCI-CNTL/PCI-LA/$1N2756 ),
    .O(\PCI-CNTL/ADX12 )
  );
  X_AND2   \PCI-CNTL/PCI-LA/$1I2708  (
    .I0(\PCI-CNTL/PCI-LA/AD7610-0000 ),
    .I1(\PCI-CNTL/PCI-LA/$1N2621 ),
    .O(\PCI-CNTL/ADX13 )
  );
  X_AND2   \PCI-CNTL/PCI-LA/$1I2705  (
    .I0(\PCI-CNTL/PCI-LA/AD7610-0000 ),
    .I1(\PCI-CNTL/PCI-LA/$1N2620 ),
    .O(\PCI-CNTL/ADX14 )
  );
  X_AND2   \PCI-CNTL/PCI-LA/$1I2701  (
    .I0(\PCI-CNTL/PCI-LA/AD7610-0000 ),
    .I1(\PCI-CNTL/PCI-LA/$1N2619 ),
    .O(\PCI-CNTL/ADX15 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LA/Q6/FDCE  (
    .CE(ADDR_VLD0),
    .CLK(CLK),
    .I(\PCI-CNTL/ADX6 ),
    .O(\PCI-CNTL/LADX6 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND4   \PCI-CNTL/PCI-LA/DEC-A/AND4  (
    .I0(\PCI-CNTL/PCI-LA/DEC-A/$1N2275 ),
    .I1(AD3),
    .I2(\PCI-CNTL/PCI-LA/DEC-A/$1N2277 ),
    .I3(AD5),
    .O(\PCI-CNTL/PCI-LA/$1N2624 )
  );
  X_INV   \PCI-CNTL/PCI-LA/DEC-A/INV2  (
    .I(AD4),
    .O(\PCI-CNTL/PCI-LA/DEC-A/$1N2277 )
  );
  X_INV   \PCI-CNTL/PCI-LA/DEC-A/INV0  (
    .I(AD2),
    .O(\PCI-CNTL/PCI-LA/DEC-A/$1N2275 )
  );
  X_AND4   \PCI-CNTL/PCI-LA/DEC-B/AND4  (
    .I0(AD2),
    .I1(AD3),
    .I2(\PCI-CNTL/PCI-LA/DEC-B/$1N2277 ),
    .I3(AD5),
    .O(\PCI-CNTL/PCI-LA/$1N2623 )
  );
  X_INV   \PCI-CNTL/PCI-LA/DEC-B/INV2  (
    .I(AD4),
    .O(\PCI-CNTL/PCI-LA/DEC-B/$1N2277 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LA/Q15/FDCE  (
    .CE(ADDR_VLD0),
    .CLK(CLK),
    .I(\PCI-CNTL/ADX15 ),
    .O(\PCI-CNTL/LADX15 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LA/Q14/FDCE  (
    .CE(ADDR_VLD0),
    .CLK(CLK),
    .I(\PCI-CNTL/ADX14 ),
    .O(\PCI-CNTL/LADX14 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LA/Q13/FDCE  (
    .CE(ADDR_VLD0),
    .CLK(CLK),
    .I(\PCI-CNTL/ADX13 ),
    .O(\PCI-CNTL/LADX13 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LA/Q12/FDCE  (
    .CE(ADDR_VLD0),
    .CLK(CLK),
    .I(\PCI-CNTL/ADX12 ),
    .O(\PCI-CNTL/LADX12 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LA/Q11/FDCE  (
    .CE(ADDR_VLD0),
    .CLK(CLK),
    .I(\PCI-CNTL/ADX11 ),
    .O(\PCI-CNTL/LADX11 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LA/Q10/FDCE  (
    .CE(ADDR_VLD0),
    .CLK(CLK),
    .I(\PCI-CNTL/ADX10 ),
    .O(\PCI-CNTL/LADX10 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LA/Q9/FDCE  (
    .CE(ADDR_VLD0),
    .CLK(CLK),
    .I(\PCI-CNTL/ADX9 ),
    .O(\PCI-CNTL/LADX9 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LA/Q8/FDCE  (
    .CE(ADDR_VLD0),
    .CLK(CLK),
    .I(\PCI-CNTL/ADX8 ),
    .O(\PCI-CNTL/LADX8 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND4   \PCI-CNTL/PCI-LA/DEC-C/AND4  (
    .I0(\PCI-CNTL/PCI-LA/DEC-C/$1N2289 ),
    .I1(\PCI-CNTL/PCI-LA/DEC-C/$1N2290 ),
    .I2(AD4),
    .I3(AD5),
    .O(\PCI-CNTL/PCI-LA/$1N2756 )
  );
  X_INV   \PCI-CNTL/PCI-LA/DEC-C/INV1  (
    .I(AD3),
    .O(\PCI-CNTL/PCI-LA/DEC-C/$1N2290 )
  );
  X_INV   \PCI-CNTL/PCI-LA/DEC-C/INV0  (
    .I(AD2),
    .O(\PCI-CNTL/PCI-LA/DEC-C/$1N2289 )
  );
  X_AND4   \PCI-CNTL/PCI-LA/DEC-F/AND4  (
    .I0(AD2),
    .I1(AD3),
    .I2(AD4),
    .I3(AD5),
    .O(\PCI-CNTL/PCI-LA/$1N2619 )
  );
  X_AND4   \PCI-CNTL/PCI-LA/DEC-D/AND4  (
    .I0(AD2),
    .I1(\PCI-CNTL/PCI-LA/DEC-D/$1N2290 ),
    .I2(AD4),
    .I3(AD5),
    .O(\PCI-CNTL/PCI-LA/$1N2621 )
  );
  X_INV   \PCI-CNTL/PCI-LA/DEC-D/INV1  (
    .I(AD3),
    .O(\PCI-CNTL/PCI-LA/DEC-D/$1N2290 )
  );
  X_AND4   \PCI-CNTL/PCI-LA/DEC-E/AND4  (
    .I0(\PCI-CNTL/PCI-LA/DEC-E/$1N2275 ),
    .I1(AD3),
    .I2(AD4),
    .I3(AD5),
    .O(\PCI-CNTL/PCI-LA/$1N2620 )
  );
  X_INV   \PCI-CNTL/PCI-LA/DEC-E/INV0  (
    .I(AD2),
    .O(\PCI-CNTL/PCI-LA/DEC-E/$1N2275 )
  );
  X_AND4   \PCI-CNTL/PCI-LA/DEC-9/AND4  (
    .I0(AD2),
    .I1(\PCI-CNTL/PCI-LA/DEC-9/$1N2276 ),
    .I2(\PCI-CNTL/PCI-LA/DEC-9/$1N2277 ),
    .I3(AD5),
    .O(\PCI-CNTL/PCI-LA/$1N2625 )
  );
  X_INV   \PCI-CNTL/PCI-LA/DEC-9/INV2  (
    .I(AD4),
    .O(\PCI-CNTL/PCI-LA/DEC-9/$1N2277 )
  );
  X_INV   \PCI-CNTL/PCI-LA/DEC-9/INV1  (
    .I(AD3),
    .O(\PCI-CNTL/PCI-LA/DEC-9/$1N2276 )
  );
  X_AND4   \PCI-CNTL/PCI-LA/DEC-8/AND4  (
    .I0(\PCI-CNTL/PCI-LA/DEC-8/$1N2275 ),
    .I1(\PCI-CNTL/PCI-LA/DEC-8/$1N2276 ),
    .I2(\PCI-CNTL/PCI-LA/DEC-8/$1N2277 ),
    .I3(AD5),
    .O(\PCI-CNTL/PCI-LA/$1N2760 )
  );
  X_INV   \PCI-CNTL/PCI-LA/DEC-8/INV2  (
    .I(AD4),
    .O(\PCI-CNTL/PCI-LA/DEC-8/$1N2277 )
  );
  X_INV   \PCI-CNTL/PCI-LA/DEC-8/INV1  (
    .I(AD3),
    .O(\PCI-CNTL/PCI-LA/DEC-8/$1N2276 )
  );
  X_INV   \PCI-CNTL/PCI-LA/DEC-8/INV0  (
    .I(AD2),
    .O(\PCI-CNTL/PCI-LA/DEC-8/$1N2275 )
  );
  X_AND4   \PCI-CNTL/PCI-LA/DEC-7/AND4  (
    .I0(AD2),
    .I1(AD3),
    .I2(AD4),
    .I3(\PCI-CNTL/PCI-LA/DEC-7/$1N2283 ),
    .O(\PCI-CNTL/PCI-LA/$1N2768 )
  );
  X_INV   \PCI-CNTL/PCI-LA/DEC-7/INV3  (
    .I(AD5),
    .O(\PCI-CNTL/PCI-LA/DEC-7/$1N2283 )
  );
  X_AND4   \PCI-CNTL/PCI-LA/DEC-6/AND4  (
    .I0(\PCI-CNTL/PCI-LA/DEC-6/$1N2275 ),
    .I1(AD3),
    .I2(AD4),
    .I3(\PCI-CNTL/PCI-LA/DEC-6/$1N2283 ),
    .O(\PCI-CNTL/PCI-LA/$1N2672 )
  );
  X_INV   \PCI-CNTL/PCI-LA/DEC-6/INV3  (
    .I(AD5),
    .O(\PCI-CNTL/PCI-LA/DEC-6/$1N2283 )
  );
  X_INV   \PCI-CNTL/PCI-LA/DEC-6/INV0  (
    .I(AD2),
    .O(\PCI-CNTL/PCI-LA/DEC-6/$1N2275 )
  );
  X_AND4   \PCI-CNTL/PCI-LA/DEC-5/AND4  (
    .I0(AD2),
    .I1(\PCI-CNTL/PCI-LA/DEC-5/$1N2276 ),
    .I2(AD4),
    .I3(\PCI-CNTL/PCI-LA/DEC-5/$1N2283 ),
    .O(\PCI-CNTL/PCI-LA/$1N2766 )
  );
  X_INV   \PCI-CNTL/PCI-LA/DEC-5/INV3  (
    .I(AD5),
    .O(\PCI-CNTL/PCI-LA/DEC-5/$1N2283 )
  );
  X_INV   \PCI-CNTL/PCI-LA/DEC-5/INV1  (
    .I(AD3),
    .O(\PCI-CNTL/PCI-LA/DEC-5/$1N2276 )
  );
  X_AND4   \PCI-CNTL/PCI-LA/DEC-4/AND4  (
    .I0(\PCI-CNTL/PCI-LA/DEC-4/$1N2275 ),
    .I1(\PCI-CNTL/PCI-LA/DEC-4/$1N2276 ),
    .I2(AD4),
    .I3(\PCI-CNTL/PCI-LA/DEC-4/$1N2283 ),
    .O(\PCI-CNTL/PCI-LA/$1N2670 )
  );
  X_INV   \PCI-CNTL/PCI-LA/DEC-4/INV3  (
    .I(AD5),
    .O(\PCI-CNTL/PCI-LA/DEC-4/$1N2283 )
  );
  X_INV   \PCI-CNTL/PCI-LA/DEC-4/INV1  (
    .I(AD3),
    .O(\PCI-CNTL/PCI-LA/DEC-4/$1N2276 )
  );
  X_INV   \PCI-CNTL/PCI-LA/DEC-4/INV0  (
    .I(AD2),
    .O(\PCI-CNTL/PCI-LA/DEC-4/$1N2275 )
  );
  X_AND4   \PCI-CNTL/PCI-LA/DEC-3/AND4  (
    .I0(AD2),
    .I1(AD3),
    .I2(\PCI-CNTL/PCI-LA/DEC-3/$1N2277 ),
    .I3(\PCI-CNTL/PCI-LA/DEC-3/$1N2283 ),
    .O(\PCI-CNTL/PCI-LA/$1N2764 )
  );
  X_INV   \PCI-CNTL/PCI-LA/DEC-3/INV3  (
    .I(AD5),
    .O(\PCI-CNTL/PCI-LA/DEC-3/$1N2283 )
  );
  X_INV   \PCI-CNTL/PCI-LA/DEC-3/INV2  (
    .I(AD4),
    .O(\PCI-CNTL/PCI-LA/DEC-3/$1N2277 )
  );
  X_AND4   \PCI-CNTL/PCI-LA/DEC-2/AND4  (
    .I0(\PCI-CNTL/PCI-LA/DEC-2/$1N2275 ),
    .I1(AD3),
    .I2(\PCI-CNTL/PCI-LA/DEC-2/$1N2277 ),
    .I3(\PCI-CNTL/PCI-LA/DEC-2/$1N2283 ),
    .O(\PCI-CNTL/PCI-LA/$1N2668 )
  );
  X_INV   \PCI-CNTL/PCI-LA/DEC-2/INV3  (
    .I(AD5),
    .O(\PCI-CNTL/PCI-LA/DEC-2/$1N2283 )
  );
  X_INV   \PCI-CNTL/PCI-LA/DEC-2/INV2  (
    .I(AD4),
    .O(\PCI-CNTL/PCI-LA/DEC-2/$1N2277 )
  );
  X_INV   \PCI-CNTL/PCI-LA/DEC-2/INV0  (
    .I(AD2),
    .O(\PCI-CNTL/PCI-LA/DEC-2/$1N2275 )
  );
  X_AND4   \PCI-CNTL/PCI-LA/DEC-0/AND4  (
    .I0(\PCI-CNTL/PCI-LA/DEC-0/$1N2275 ),
    .I1(\PCI-CNTL/PCI-LA/DEC-0/$1N2276 ),
    .I2(\PCI-CNTL/PCI-LA/DEC-0/$1N2277 ),
    .I3(\PCI-CNTL/PCI-LA/DEC-0/$1N2283 ),
    .O(\PCI-CNTL/PCI-LA/$1N2666 )
  );
  X_INV   \PCI-CNTL/PCI-LA/DEC-0/INV3  (
    .I(AD5),
    .O(\PCI-CNTL/PCI-LA/DEC-0/$1N2283 )
  );
  X_INV   \PCI-CNTL/PCI-LA/DEC-0/INV2  (
    .I(AD4),
    .O(\PCI-CNTL/PCI-LA/DEC-0/$1N2277 )
  );
  X_INV   \PCI-CNTL/PCI-LA/DEC-0/INV1  (
    .I(AD3),
    .O(\PCI-CNTL/PCI-LA/DEC-0/$1N2276 )
  );
  X_INV   \PCI-CNTL/PCI-LA/DEC-0/INV0  (
    .I(AD2),
    .O(\PCI-CNTL/PCI-LA/DEC-0/$1N2275 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LA/Q2/FDCE  (
    .CE(ADDR_VLD0),
    .CLK(CLK),
    .I(\PCI-CNTL/ADX2 ),
    .O(\PCI-CNTL/LADX2 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LA/Q3/FDCE  (
    .CE(ADDR_VLD0),
    .CLK(CLK),
    .I(\PCI-CNTL/ADX3 ),
    .O(\PCI-CNTL/LADX3 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LA/Q1/FDCE  (
    .CE(ADDR_VLD0),
    .CLK(CLK),
    .I(\PCI-CNTL/ADX1 ),
    .O(\PCI-CNTL/LADX1 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LA/Q0/FDCE  (
    .CE(ADDR_VLD0),
    .CLK(CLK),
    .I(\PCI-CNTL/ADX0 ),
    .O(\PCI-CNTL/LADX0 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_INV   \PCI-CNTL/PCI-LA/DEC-1/INV1  (
    .I(AD3),
    .O(\PCI-CNTL/PCI-LA/DEC-1/$1N2280 )
  );
  X_INV   \PCI-CNTL/PCI-LA/DEC-1/INV2  (
    .I(AD4),
    .O(\PCI-CNTL/PCI-LA/DEC-1/$1N2278 )
  );
  X_INV   \PCI-CNTL/PCI-LA/DEC-1/INV3  (
    .I(AD5),
    .O(\PCI-CNTL/PCI-LA/DEC-1/$1N2277 )
  );
  X_AND4   \PCI-CNTL/PCI-LA/DEC-1/AND4  (
    .I0(AD2),
    .I1(\PCI-CNTL/PCI-LA/DEC-1/$1N2280 ),
    .I2(\PCI-CNTL/PCI-LA/DEC-1/$1N2278 ),
    .I3(\PCI-CNTL/PCI-LA/DEC-1/$1N2277 ),
    .O(\PCI-CNTL/PCI-LA/$1N2762 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LA/Q4/FDCE  (
    .CE(ADDR_VLD0),
    .CLK(CLK),
    .I(\PCI-CNTL/ADX4 ),
    .O(\PCI-CNTL/LADX4 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LA/Q5/FDCE  (
    .CE(ADDR_VLD0),
    .CLK(CLK),
    .I(\PCI-CNTL/ADX5 ),
    .O(\PCI-CNTL/LADX5 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LA/Q7/FDCE  (
    .CE(ADDR_VLD0),
    .CLK(CLK),
    .I(\PCI-CNTL/ADX7 ),
    .O(\PCI-CNTL/LADX7 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND4   \PCI-CNTL/PCI-LA/0000/AND4  (
    .I0(\PCI-CNTL/PCI-LA/0000/$1N2275 ),
    .I1(\PCI-CNTL/PCI-LA/0000/$1N2276 ),
    .I2(\PCI-CNTL/PCI-LA/0000/$1N2277 ),
    .I3(\PCI-CNTL/PCI-LA/0000/$1N2283 ),
    .O(\PCI-CNTL/PCI-LA/AD7610-0000 )
  );
  X_INV   \PCI-CNTL/PCI-LA/0000/INV3  (
    .I(AD7),
    .O(\PCI-CNTL/PCI-LA/0000/$1N2283 )
  );
  X_INV   \PCI-CNTL/PCI-LA/0000/INV2  (
    .I(AD6),
    .O(\PCI-CNTL/PCI-LA/0000/$1N2277 )
  );
  X_INV   \PCI-CNTL/PCI-LA/0000/INV1  (
    .I(AD1),
    .O(\PCI-CNTL/PCI-LA/0000/$1N2276 )
  );
  X_INV   \PCI-CNTL/PCI-LA/0000/INV0  (
    .I(AD0),
    .O(\PCI-CNTL/PCI-LA/0000/$1N2275 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LA/LA4/FDCE  (
    .CE(ADDR_VLD0),
    .CLK(CLK),
    .I(AD4),
    .O(NlwRenamedSig_OI_ADDR4),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LA/LA5/FDCE  (
    .CE(ADDR_VLD0),
    .CLK(CLK),
    .I(AD5),
    .O(NlwRenamedSig_OI_ADDR5),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LA/LA3/FDCE  (
    .CE(ADDR_VLD0),
    .CLK(CLK),
    .I(AD3),
    .O(NlwRenamedSig_OI_ADDR3),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LA/LA2/FDCE  (
    .CE(ADDR_VLD0),
    .CLK(CLK),
    .I(AD2),
    .O(NlwRenamedSig_OI_ADDR2),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LA/LA1/FDCE  (
    .CE(ADDR_VLD0),
    .CLK(CLK),
    .I(AD1),
    .O(NlwRenamedSig_OI_ADDR1),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LA/LA0/FDCE  (
    .CE(ADDR_VLD0),
    .CLK(CLK),
    .I(AD0),
    .O(NlwRenamedSig_OI_ADDR0),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LA/LA6/FDCE  (
    .CE(ADDR_VLD0),
    .CLK(CLK),
    .I(AD6),
    .O(NlwRenamedSig_OI_ADDR6),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LA/LA7/FDCE  (
    .CE(ADDR_VLD0),
    .CLK(CLK),
    .I(AD7),
    .O(NlwRenamedSig_OI_ADDR7),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LA/LA8/FDCE  (
    .CE(ADDR_VLD0),
    .CLK(CLK),
    .I(AD8),
    .O(NlwRenamedSig_OI_ADDR8),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LA/LA15/FDCE  (
    .CE(ADDR_VLD0),
    .CLK(CLK),
    .I(AD15),
    .O(NlwRenamedSig_OI_ADDR15),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LA/LA14/FDCE  (
    .CE(ADDR_VLD0),
    .CLK(CLK),
    .I(AD14),
    .O(NlwRenamedSig_OI_ADDR14),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LA/LA13/FDCE  (
    .CE(ADDR_VLD0),
    .CLK(CLK),
    .I(AD13),
    .O(NlwRenamedSig_OI_ADDR13),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LA/LA9/FDCE  (
    .CE(ADDR_VLD0),
    .CLK(CLK),
    .I(AD9),
    .O(NlwRenamedSig_OI_ADDR9),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LA/LA10/FDCE  (
    .CE(ADDR_VLD0),
    .CLK(CLK),
    .I(AD10),
    .O(NlwRenamedSig_OI_ADDR10),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LA/LA11/FDCE  (
    .CE(ADDR_VLD0),
    .CLK(CLK),
    .I(AD11),
    .O(NlwRenamedSig_OI_ADDR11),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LA/LA12/FDCE  (
    .CE(ADDR_VLD0),
    .CLK(CLK),
    .I(AD12),
    .O(NlwRenamedSig_OI_ADDR12),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LA/LA20/FDCE  (
    .CE(ADDR_VLD0),
    .CLK(CLK),
    .I(AD20),
    .O(NlwRenamedSig_OI_ADDR20),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LA/LA19/FDCE  (
    .CE(ADDR_VLD0),
    .CLK(CLK),
    .I(AD19),
    .O(NlwRenamedSig_OI_ADDR19),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LA/LA18/FDCE  (
    .CE(ADDR_VLD0),
    .CLK(CLK),
    .I(AD18),
    .O(NlwRenamedSig_OI_ADDR18),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LA/LA21/FDCE  (
    .CE(ADDR_VLD0),
    .CLK(CLK),
    .I(AD21),
    .O(NlwRenamedSig_OI_ADDR21),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LA/LA22/FDCE  (
    .CE(ADDR_VLD0),
    .CLK(CLK),
    .I(AD22),
    .O(NlwRenamedSig_OI_ADDR22),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LA/LA23/FDCE  (
    .CE(ADDR_VLD0),
    .CLK(CLK),
    .I(AD23),
    .O(NlwRenamedSig_OI_ADDR23),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LA/LA16/FDCE  (
    .CE(ADDR_VLD0),
    .CLK(CLK),
    .I(AD16),
    .O(NlwRenamedSig_OI_ADDR16),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LA/LA17/FDCE  (
    .CE(ADDR_VLD0),
    .CLK(CLK),
    .I(AD17),
    .O(NlwRenamedSig_OI_ADDR17),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LA/LA31/FDCE  (
    .CE(ADDR_VLD0),
    .CLK(CLK),
    .I(AD31),
    .O(NlwRenamedSig_OI_ADDR31),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LA/LA30/FDCE  (
    .CE(ADDR_VLD0),
    .CLK(CLK),
    .I(AD30),
    .O(NlwRenamedSig_OI_ADDR30),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LA/LA29/FDCE  (
    .CE(ADDR_VLD0),
    .CLK(CLK),
    .I(AD29),
    .O(NlwRenamedSig_OI_ADDR29),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LA/LA26/FDCE  (
    .CE(ADDR_VLD0),
    .CLK(CLK),
    .I(AD26),
    .O(NlwRenamedSig_OI_ADDR26),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LA/LA27/FDCE  (
    .CE(ADDR_VLD0),
    .CLK(CLK),
    .I(AD27),
    .O(NlwRenamedSig_OI_ADDR27),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LA/LA28/FDCE  (
    .CE(ADDR_VLD0),
    .CLK(CLK),
    .I(AD28),
    .O(NlwRenamedSig_OI_ADDR28),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LA/LA25/FDCE  (
    .CE(ADDR_VLD0),
    .CLK(CLK),
    .I(AD25),
    .O(NlwRenamedSig_OI_ADDR25),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LA/LA24/FDCE  (
    .CE(ADDR_VLD0),
    .CLK(CLK),
    .I(AD24),
    .O(NlwRenamedSig_OI_ADDR24),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LC/CFG_CYC  (
    .CE(VCC),
    .CLK(CLK),
    .I(\PCI-CNTL/PCI-LC/NS_CFG_CYC ),
    .O(\PCI-CNTL/CFG_CYC ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND2   \PCI-CNTL/PCI-LC/$2I3221  (
    .I0(ADDR_VLD1),
    .I1(\PCI-CNTL/PCI-LC/$2N3210 ),
    .O(\PCI-CNTL/NS_CFG_HIT )
  );
  X_AND2   \PCI-CNTL/PCI-LC/$2I3214  (
    .I0(\PCI-CNTL/PCI-LC/$2N3209 ),
    .I1(\PCI-CNTL/PCI-LC/RW_CFG ),
    .O(\PCI-CNTL/PCI-LC/$2N3210 )
  );
  X_AND2   \PCI-CNTL/PCI-LC/$2I3213  (
    .I0(IDSEL),
    .I1(\PCI-CNTL/PCI-LC/TYPE00 ),
    .O(\PCI-CNTL/PCI-LC/$2N3209 )
  );
  X_AND2   \PCI-CNTL/PCI-LC/$2I3201  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-LC/$2I3201/I0 ),
    .I1(\NlwInverterSignal_PCI-CNTL/PCI-LC/$2I3201/I1 ),
    .O(\PCI-CNTL/PCI-LC/TYPE00 )
  );
  X_AND3   \PCI-CNTL/PCI-LC/$2I3192  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-LC/$2I3192/I0 ),
    .I1(CBE_IN1),
    .I2(CBE_IN3),
    .O(\PCI-CNTL/PCI-LC/RW_CFG )
  );
  X_AND2   \PCI-CNTL/PCI-LC/$2I3076  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-LC/$2I3076/I0 ),
    .I1(\PCI-CNTL/CFG_CYC ),
    .O(\PCI-CNTL/PCI-LC/$2N2912 )
  );
  X_OR2   \PCI-CNTL/PCI-LC/$2I3073  (
    .I0(\PCI-CNTL/NS_CFG_HIT ),
    .I1(\PCI-CNTL/PCI-LC/$2N2912 ),
    .O(\PCI-CNTL/PCI-LC/NS_CFG_CYC )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LC/CFG_HIT  (
    .CE(VCC),
    .CLK(CLK),
    .I(\PCI-CNTL/NS_CFG_HIT ),
    .O(NlwRenamedSig_OI_CFG_HIT),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LC/Q6/FDCE  (
    .CE(ADDR_VLD1),
    .CLK(CLK),
    .I(\PCI-CNTL/CMD6 ),
    .O(NlwRenamedSig_OI_PCI_CMD6),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LC/Q7/FDCE  (
    .CE(ADDR_VLD1),
    .CLK(CLK),
    .I(\PCI-CNTL/CMD7 ),
    .O(NlwRenamedSig_OI_PCI_CMD7),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LC/Q5/FDCE  (
    .CE(ADDR_VLD1),
    .CLK(CLK),
    .I(\PCI-CNTL/CMD5 ),
    .O(NlwRenamedSig_OI_PCI_CMD5),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LC/Q4/FDCE  (
    .CE(ADDR_VLD1),
    .CLK(CLK),
    .I(\PCI-CNTL/CMD4 ),
    .O(NlwRenamedSig_OI_PCI_CMD4),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LC/Q2/FDCE  (
    .CE(ADDR_VLD1),
    .CLK(CLK),
    .I(\PCI-CNTL/CMD2 ),
    .O(NlwRenamedSig_OI_PCI_CMD2),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LC/Q3/FDCE  (
    .CE(ADDR_VLD1),
    .CLK(CLK),
    .I(\PCI-CNTL/CMD3 ),
    .O(NlwRenamedSig_OI_PCI_CMD3),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LC/Q1/FDCE  (
    .CE(ADDR_VLD1),
    .CLK(CLK),
    .I(\PCI-CNTL/CMD1 ),
    .O(NlwRenamedSig_OI_PCI_CMD1),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LC/Q0/FDCE  (
    .CE(ADDR_VLD1),
    .CLK(CLK),
    .I(\PCI-CNTL/CMD0 ),
    .O(NlwRenamedSig_OI_PCI_CMD0),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND4   \PCI-CNTL/PCI-LC/DEC-E/AND4  (
    .I0(\PCI-CNTL/PCI-LC/DEC-E/$1N2275 ),
    .I1(CBE_IN1),
    .I2(CBE_IN2),
    .I3(CBE_IN3),
    .O(\PCI-CNTL/CMD14 )
  );
  X_INV   \PCI-CNTL/PCI-LC/DEC-E/INV0  (
    .I(CBE_IN0),
    .O(\PCI-CNTL/PCI-LC/DEC-E/$1N2275 )
  );
  X_AND4   \PCI-CNTL/PCI-LC/DEC-D/AND4  (
    .I0(CBE_IN0),
    .I1(\PCI-CNTL/PCI-LC/DEC-D/$1N2290 ),
    .I2(CBE_IN2),
    .I3(CBE_IN3),
    .O(\PCI-CNTL/CMD13 )
  );
  X_INV   \PCI-CNTL/PCI-LC/DEC-D/INV1  (
    .I(CBE_IN1),
    .O(\PCI-CNTL/PCI-LC/DEC-D/$1N2290 )
  );
  X_AND4   \PCI-CNTL/PCI-LC/DEC-F/AND4  (
    .I0(CBE_IN0),
    .I1(CBE_IN1),
    .I2(CBE_IN2),
    .I3(CBE_IN3),
    .O(\PCI-CNTL/CMD15 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LC/Q12/FDCE  (
    .CE(ADDR_VLD1),
    .CLK(CLK),
    .I(\PCI-CNTL/CMD12 ),
    .O(NlwRenamedSig_OI_PCI_CMD12),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LC/Q13/FDCE  (
    .CE(ADDR_VLD1),
    .CLK(CLK),
    .I(\PCI-CNTL/CMD13 ),
    .O(NlwRenamedSig_OI_PCI_CMD13),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LC/Q15/FDCE  (
    .CE(ADDR_VLD1),
    .CLK(CLK),
    .I(\PCI-CNTL/CMD15 ),
    .O(NlwRenamedSig_OI_PCI_CMD15),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LC/Q14/FDCE  (
    .CE(ADDR_VLD1),
    .CLK(CLK),
    .I(\PCI-CNTL/CMD14 ),
    .O(NlwRenamedSig_OI_PCI_CMD14),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND4   \PCI-CNTL/PCI-LC/DEC-C/AND4  (
    .I0(\PCI-CNTL/PCI-LC/DEC-C/$1N2289 ),
    .I1(\PCI-CNTL/PCI-LC/DEC-C/$1N2290 ),
    .I2(CBE_IN2),
    .I3(CBE_IN3),
    .O(\PCI-CNTL/CMD12 )
  );
  X_INV   \PCI-CNTL/PCI-LC/DEC-C/INV1  (
    .I(CBE_IN1),
    .O(\PCI-CNTL/PCI-LC/DEC-C/$1N2290 )
  );
  X_INV   \PCI-CNTL/PCI-LC/DEC-C/INV0  (
    .I(CBE_IN0),
    .O(\PCI-CNTL/PCI-LC/DEC-C/$1N2289 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LC/Q8/FDCE  (
    .CE(ADDR_VLD1),
    .CLK(CLK),
    .I(\PCI-CNTL/CMD8 ),
    .O(NlwRenamedSig_OI_PCI_CMD8),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LC/Q9/FDCE  (
    .CE(ADDR_VLD1),
    .CLK(CLK),
    .I(\PCI-CNTL/CMD9 ),
    .O(NlwRenamedSig_OI_PCI_CMD9),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LC/Q11/FDCE  (
    .CE(ADDR_VLD1),
    .CLK(CLK),
    .I(\PCI-CNTL/CMD11 ),
    .O(NlwRenamedSig_OI_PCI_CMD11),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LC/Q10/FDCE  (
    .CE(ADDR_VLD1),
    .CLK(CLK),
    .I(\PCI-CNTL/CMD10 ),
    .O(NlwRenamedSig_OI_PCI_CMD10),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND4   \PCI-CNTL/PCI-LC/DEC-0/AND4  (
    .I0(\PCI-CNTL/PCI-LC/DEC-0/$1N2275 ),
    .I1(\PCI-CNTL/PCI-LC/DEC-0/$1N2276 ),
    .I2(\PCI-CNTL/PCI-LC/DEC-0/$1N2277 ),
    .I3(\PCI-CNTL/PCI-LC/DEC-0/$1N2283 ),
    .O(\PCI-CNTL/CMD0 )
  );
  X_INV   \PCI-CNTL/PCI-LC/DEC-0/INV3  (
    .I(CBE_IN3),
    .O(\PCI-CNTL/PCI-LC/DEC-0/$1N2283 )
  );
  X_INV   \PCI-CNTL/PCI-LC/DEC-0/INV2  (
    .I(CBE_IN2),
    .O(\PCI-CNTL/PCI-LC/DEC-0/$1N2277 )
  );
  X_INV   \PCI-CNTL/PCI-LC/DEC-0/INV1  (
    .I(CBE_IN1),
    .O(\PCI-CNTL/PCI-LC/DEC-0/$1N2276 )
  );
  X_INV   \PCI-CNTL/PCI-LC/DEC-0/INV0  (
    .I(CBE_IN0),
    .O(\PCI-CNTL/PCI-LC/DEC-0/$1N2275 )
  );
  X_INV   \PCI-CNTL/PCI-LC/DEC-1/INV1  (
    .I(CBE_IN1),
    .O(\PCI-CNTL/PCI-LC/DEC-1/$1N2280 )
  );
  X_INV   \PCI-CNTL/PCI-LC/DEC-1/INV2  (
    .I(CBE_IN2),
    .O(\PCI-CNTL/PCI-LC/DEC-1/$1N2278 )
  );
  X_INV   \PCI-CNTL/PCI-LC/DEC-1/INV3  (
    .I(CBE_IN3),
    .O(\PCI-CNTL/PCI-LC/DEC-1/$1N2277 )
  );
  X_AND4   \PCI-CNTL/PCI-LC/DEC-1/AND4  (
    .I0(CBE_IN0),
    .I1(\PCI-CNTL/PCI-LC/DEC-1/$1N2280 ),
    .I2(\PCI-CNTL/PCI-LC/DEC-1/$1N2278 ),
    .I3(\PCI-CNTL/PCI-LC/DEC-1/$1N2277 ),
    .O(\PCI-CNTL/CMD1 )
  );
  X_AND4   \PCI-CNTL/PCI-LC/DEC-2/AND4  (
    .I0(\PCI-CNTL/PCI-LC/DEC-2/$1N2275 ),
    .I1(CBE_IN1),
    .I2(\PCI-CNTL/PCI-LC/DEC-2/$1N2277 ),
    .I3(\PCI-CNTL/PCI-LC/DEC-2/$1N2283 ),
    .O(\PCI-CNTL/CMD2 )
  );
  X_INV   \PCI-CNTL/PCI-LC/DEC-2/INV3  (
    .I(CBE_IN3),
    .O(\PCI-CNTL/PCI-LC/DEC-2/$1N2283 )
  );
  X_INV   \PCI-CNTL/PCI-LC/DEC-2/INV2  (
    .I(CBE_IN2),
    .O(\PCI-CNTL/PCI-LC/DEC-2/$1N2277 )
  );
  X_INV   \PCI-CNTL/PCI-LC/DEC-2/INV0  (
    .I(CBE_IN0),
    .O(\PCI-CNTL/PCI-LC/DEC-2/$1N2275 )
  );
  X_AND4   \PCI-CNTL/PCI-LC/DEC-3/AND4  (
    .I0(CBE_IN0),
    .I1(CBE_IN1),
    .I2(\PCI-CNTL/PCI-LC/DEC-3/$1N2277 ),
    .I3(\PCI-CNTL/PCI-LC/DEC-3/$1N2283 ),
    .O(\PCI-CNTL/CMD3 )
  );
  X_INV   \PCI-CNTL/PCI-LC/DEC-3/INV3  (
    .I(CBE_IN3),
    .O(\PCI-CNTL/PCI-LC/DEC-3/$1N2283 )
  );
  X_INV   \PCI-CNTL/PCI-LC/DEC-3/INV2  (
    .I(CBE_IN2),
    .O(\PCI-CNTL/PCI-LC/DEC-3/$1N2277 )
  );
  X_AND4   \PCI-CNTL/PCI-LC/DEC-4/AND4  (
    .I0(\PCI-CNTL/PCI-LC/DEC-4/$1N2275 ),
    .I1(\PCI-CNTL/PCI-LC/DEC-4/$1N2276 ),
    .I2(CBE_IN2),
    .I3(\PCI-CNTL/PCI-LC/DEC-4/$1N2283 ),
    .O(\PCI-CNTL/CMD4 )
  );
  X_INV   \PCI-CNTL/PCI-LC/DEC-4/INV3  (
    .I(CBE_IN3),
    .O(\PCI-CNTL/PCI-LC/DEC-4/$1N2283 )
  );
  X_INV   \PCI-CNTL/PCI-LC/DEC-4/INV1  (
    .I(CBE_IN1),
    .O(\PCI-CNTL/PCI-LC/DEC-4/$1N2276 )
  );
  X_INV   \PCI-CNTL/PCI-LC/DEC-4/INV0  (
    .I(CBE_IN0),
    .O(\PCI-CNTL/PCI-LC/DEC-4/$1N2275 )
  );
  X_AND4   \PCI-CNTL/PCI-LC/DEC-5/AND4  (
    .I0(CBE_IN0),
    .I1(\PCI-CNTL/PCI-LC/DEC-5/$1N2276 ),
    .I2(CBE_IN2),
    .I3(\PCI-CNTL/PCI-LC/DEC-5/$1N2283 ),
    .O(\PCI-CNTL/CMD5 )
  );
  X_INV   \PCI-CNTL/PCI-LC/DEC-5/INV3  (
    .I(CBE_IN3),
    .O(\PCI-CNTL/PCI-LC/DEC-5/$1N2283 )
  );
  X_INV   \PCI-CNTL/PCI-LC/DEC-5/INV1  (
    .I(CBE_IN1),
    .O(\PCI-CNTL/PCI-LC/DEC-5/$1N2276 )
  );
  X_AND4   \PCI-CNTL/PCI-LC/DEC-6/AND4  (
    .I0(\PCI-CNTL/PCI-LC/DEC-6/$1N2275 ),
    .I1(CBE_IN1),
    .I2(CBE_IN2),
    .I3(\PCI-CNTL/PCI-LC/DEC-6/$1N2283 ),
    .O(\PCI-CNTL/CMD6 )
  );
  X_INV   \PCI-CNTL/PCI-LC/DEC-6/INV3  (
    .I(CBE_IN3),
    .O(\PCI-CNTL/PCI-LC/DEC-6/$1N2283 )
  );
  X_INV   \PCI-CNTL/PCI-LC/DEC-6/INV0  (
    .I(CBE_IN0),
    .O(\PCI-CNTL/PCI-LC/DEC-6/$1N2275 )
  );
  X_AND4   \PCI-CNTL/PCI-LC/DEC-7/AND4  (
    .I0(CBE_IN0),
    .I1(CBE_IN1),
    .I2(CBE_IN2),
    .I3(\PCI-CNTL/PCI-LC/DEC-7/$1N2283 ),
    .O(\PCI-CNTL/CMD7 )
  );
  X_INV   \PCI-CNTL/PCI-LC/DEC-7/INV3  (
    .I(CBE_IN3),
    .O(\PCI-CNTL/PCI-LC/DEC-7/$1N2283 )
  );
  X_AND4   \PCI-CNTL/PCI-LC/DEC-8/AND4  (
    .I0(\PCI-CNTL/PCI-LC/DEC-8/$1N2275 ),
    .I1(\PCI-CNTL/PCI-LC/DEC-8/$1N2276 ),
    .I2(\PCI-CNTL/PCI-LC/DEC-8/$1N2277 ),
    .I3(CBE_IN3),
    .O(\PCI-CNTL/CMD8 )
  );
  X_INV   \PCI-CNTL/PCI-LC/DEC-8/INV2  (
    .I(CBE_IN2),
    .O(\PCI-CNTL/PCI-LC/DEC-8/$1N2277 )
  );
  X_INV   \PCI-CNTL/PCI-LC/DEC-8/INV1  (
    .I(CBE_IN1),
    .O(\PCI-CNTL/PCI-LC/DEC-8/$1N2276 )
  );
  X_INV   \PCI-CNTL/PCI-LC/DEC-8/INV0  (
    .I(CBE_IN0),
    .O(\PCI-CNTL/PCI-LC/DEC-8/$1N2275 )
  );
  X_AND4   \PCI-CNTL/PCI-LC/DEC-9/AND4  (
    .I0(CBE_IN0),
    .I1(\PCI-CNTL/PCI-LC/DEC-9/$1N2276 ),
    .I2(\PCI-CNTL/PCI-LC/DEC-9/$1N2277 ),
    .I3(CBE_IN3),
    .O(\PCI-CNTL/CMD9 )
  );
  X_INV   \PCI-CNTL/PCI-LC/DEC-9/INV2  (
    .I(CBE_IN2),
    .O(\PCI-CNTL/PCI-LC/DEC-9/$1N2277 )
  );
  X_INV   \PCI-CNTL/PCI-LC/DEC-9/INV1  (
    .I(CBE_IN1),
    .O(\PCI-CNTL/PCI-LC/DEC-9/$1N2276 )
  );
  X_AND4   \PCI-CNTL/PCI-LC/DEC-A/AND4  (
    .I0(\PCI-CNTL/PCI-LC/DEC-A/$1N2275 ),
    .I1(CBE_IN1),
    .I2(\PCI-CNTL/PCI-LC/DEC-A/$1N2277 ),
    .I3(CBE_IN3),
    .O(\PCI-CNTL/CMD10 )
  );
  X_INV   \PCI-CNTL/PCI-LC/DEC-A/INV2  (
    .I(CBE_IN2),
    .O(\PCI-CNTL/PCI-LC/DEC-A/$1N2277 )
  );
  X_INV   \PCI-CNTL/PCI-LC/DEC-A/INV0  (
    .I(CBE_IN0),
    .O(\PCI-CNTL/PCI-LC/DEC-A/$1N2275 )
  );
  X_AND4   \PCI-CNTL/PCI-LC/DEC-B/AND4  (
    .I0(CBE_IN0),
    .I1(CBE_IN1),
    .I2(\PCI-CNTL/PCI-LC/DEC-B/$1N2277 ),
    .I3(CBE_IN3),
    .O(\PCI-CNTL/CMD11 )
  );
  X_INV   \PCI-CNTL/PCI-LC/DEC-B/INV2  (
    .I(CBE_IN2),
    .O(\PCI-CNTL/PCI-LC/DEC-B/$1N2277 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LC/LC0/FDCE  (
    .CE(ADDR_VLD1),
    .CLK(CLK),
    .I(CBE_IN0),
    .O(NlwRenamedSig_OI_S_WRDN),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-LC/LC1/FDCE  (
    .CE(ADDR_VLD1),
    .CLK(CLK),
    .I(CBE_IN0),
    .O(S_WRDN_DUP),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND2   \PCI-CNTL/PCI-OE/$2I940  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OE/$2I940/I0 ),
    .I1(\PCI-CNTL/PCI-OE/$2N942 ),
    .O(\PCI-CNTL/PCI-OE/UCS )
  );
  X_AND2   \PCI-CNTL/PCI-OE/$2I934  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OE/$2I934/I0 ),
    .I1(\PCI-CNTL/PCI-OE/10H ),
    .O(\PCI-CNTL/PCI-OE/$2N755 )
  );
  X_AND2   \PCI-CNTL/PCI-OE/$2I933  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OE/$2I933/I0 ),
    .I1(\PCI-CNTL/PCI-OE/14H ),
    .O(\PCI-CNTL/PCI-OE/$2N754 )
  );
  X_AND2   \PCI-CNTL/PCI-OE/$2I932  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OE/$2I932/I0 ),
    .I1(\PCI-CNTL/PCI-OE/18H ),
    .O(\PCI-CNTL/PCI-OE/$2N753 )
  );
  X_OR2   \PCI-CNTL/PCI-OE/$2I790  (
    .I0(\PCI-CNTL/PCI-OE/$2N791 ),
    .I1(\PCI-CNTL/PCI-OE/UCS ),
    .O(\PCI-CNTL/PCI-OE/$2N795 )
  );
  X_AND2   \PCI-CNTL/PCI-OE/$2I788  (
    .I0(\PCI-CNTL/PCI-OE/LCS ),
    .I1(\PCI-CNTL/PCI-OE/X ),
    .O(\PCI-CNTL/PCI-OE/$2N791 )
  );
  X_AND2   \PCI-CNTL/PCI-OE/$2I777  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OE/$2I777/I0 ),
    .I1(\NlwInverterSignal_PCI-CNTL/PCI-OE/$2I777/I1 ),
    .O(\PCI-CNTL/PCI-OE/LCS )
  );
  X_OR2   \PCI-CNTL/PCI-OE/$2I766  (
    .I0(NlwRenamedSig_OI_ADDR6),
    .I1(NlwRenamedSig_OI_ADDR7),
    .O(\PCI-CNTL/PCI-OE/$2N942 )
  );
  X_AND4   \PCI-CNTL/PCI-OE/$2I592  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OE/$2I592/I0 ),
    .I1(NlwRenamedSig_OI_CFG_HIT),
    .I2(NlwRenamedSig_OI_PCI_CMD10),
    .I3(\PCI-CNTL/PCI-OE/$2N795 ),
    .O(\PCI-CNTL/PCI-OE/NS_OE_ROM )
  );
  X_BUF   \PCI-CNTL/PCI-OE/OE15/$1I320  (
    .I(\PCI-CNTL/PCI-OE/OE15/Q ),
    .O(OE15)
  );
  X_BUF   \PCI-CNTL/PCI-OE/OE15/$1I311  (
    .I(\PCI-CNTL/END ),
    .O(\PCI-CNTL/PCI-OE/OE15/S )
  );
  X_BUF   \PCI-CNTL/PCI-OE/OE15/$1I310  (
    .I(\PCI-CNTL/PCI-OE/OE15/NS_OE ),
    .O(\PCI-CNTL/PCI-OE/OE15/R )
  );
  X_BUF   \PCI-CNTL/PCI-OE/OE15/$1I309  (
    .I(CLK),
    .O(\PCI-CNTL/PCI-OE/OE15/C )
  );
  X_AND2   \PCI-CNTL/PCI-OE/OE15/$1I307  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OE/OE15/$1I307/I0 ),
    .I1(\PCI-CNTL/PCI-OE/OE15/Q ),
    .O(\PCI-CNTL/PCI-OE/OE15/$1N301 )
  );
  X_OR2   \PCI-CNTL/PCI-OE/OE15/$1I306  (
    .I0(\PCI-CNTL/PCI-OE/OE15/S ),
    .I1(\PCI-CNTL/PCI-OE/OE15/$1N301 ),
    .O(\PCI-CNTL/PCI-OE/OE15/D )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-CNTL/PCI-OE/OE15/FDPE  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(\PCI-CNTL/PCI-OE/OE15/C ),
    .I(\PCI-CNTL/PCI-OE/OE15/D ),
    .O(\PCI-CNTL/PCI-OE/OE15/Q ),
    .RST(GND)
  );
  X_AND4   \PCI-CNTL/PCI-OE/OE15/$1I296  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OE/OE15/$1I296/I0 ),
    .I1(NlwRenamedSig_OI_PCI_CMD10),
    .I2(\PCI-CNTL/LADX15 ),
    .I3(NlwRenamedSig_OI_CFG_HIT),
    .O(\PCI-CNTL/PCI-OE/OE15/NS_OE )
  );
  X_BUF   \PCI-CNTL/PCI-OE/OE7/$1I320  (
    .I(\PCI-CNTL/PCI-OE/OE7/Q ),
    .O(OE7)
  );
  X_BUF   \PCI-CNTL/PCI-OE/OE7/$1I311  (
    .I(\PCI-CNTL/END ),
    .O(\PCI-CNTL/PCI-OE/OE7/S )
  );
  X_BUF   \PCI-CNTL/PCI-OE/OE7/$1I310  (
    .I(\PCI-CNTL/PCI-OE/OE7/NS_OE ),
    .O(\PCI-CNTL/PCI-OE/OE7/R )
  );
  X_BUF   \PCI-CNTL/PCI-OE/OE7/$1I309  (
    .I(CLK),
    .O(\PCI-CNTL/PCI-OE/OE7/C )
  );
  X_AND2   \PCI-CNTL/PCI-OE/OE7/$1I307  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OE/OE7/$1I307/I0 ),
    .I1(\PCI-CNTL/PCI-OE/OE7/Q ),
    .O(\PCI-CNTL/PCI-OE/OE7/$1N301 )
  );
  X_OR2   \PCI-CNTL/PCI-OE/OE7/$1I306  (
    .I0(\PCI-CNTL/PCI-OE/OE7/S ),
    .I1(\PCI-CNTL/PCI-OE/OE7/$1N301 ),
    .O(\PCI-CNTL/PCI-OE/OE7/D )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-CNTL/PCI-OE/OE7/FDPE  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(\PCI-CNTL/PCI-OE/OE7/C ),
    .I(\PCI-CNTL/PCI-OE/OE7/D ),
    .O(\PCI-CNTL/PCI-OE/OE7/Q ),
    .RST(GND)
  );
  X_AND4   \PCI-CNTL/PCI-OE/OE7/$1I296  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OE/OE7/$1I296/I0 ),
    .I1(NlwRenamedSig_OI_PCI_CMD10),
    .I2(\PCI-CNTL/LADX7 ),
    .I3(NlwRenamedSig_OI_CFG_HIT),
    .O(\PCI-CNTL/PCI-OE/OE7/NS_OE )
  );
  X_BUF   \PCI-CNTL/PCI-OE/OE6/$1I320  (
    .I(\PCI-CNTL/PCI-OE/OE6/Q ),
    .O(OE6)
  );
  X_BUF   \PCI-CNTL/PCI-OE/OE6/$1I311  (
    .I(\PCI-CNTL/END ),
    .O(\PCI-CNTL/PCI-OE/OE6/S )
  );
  X_BUF   \PCI-CNTL/PCI-OE/OE6/$1I310  (
    .I(\PCI-CNTL/PCI-OE/OE6/NS_OE ),
    .O(\PCI-CNTL/PCI-OE/OE6/R )
  );
  X_BUF   \PCI-CNTL/PCI-OE/OE6/$1I309  (
    .I(CLK),
    .O(\PCI-CNTL/PCI-OE/OE6/C )
  );
  X_AND2   \PCI-CNTL/PCI-OE/OE6/$1I307  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OE/OE6/$1I307/I0 ),
    .I1(\PCI-CNTL/PCI-OE/OE6/Q ),
    .O(\PCI-CNTL/PCI-OE/OE6/$1N301 )
  );
  X_OR2   \PCI-CNTL/PCI-OE/OE6/$1I306  (
    .I0(\PCI-CNTL/PCI-OE/OE6/S ),
    .I1(\PCI-CNTL/PCI-OE/OE6/$1N301 ),
    .O(\PCI-CNTL/PCI-OE/OE6/D )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-CNTL/PCI-OE/OE6/FDPE  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(\PCI-CNTL/PCI-OE/OE6/C ),
    .I(\PCI-CNTL/PCI-OE/OE6/D ),
    .O(\PCI-CNTL/PCI-OE/OE6/Q ),
    .RST(GND)
  );
  X_AND4   \PCI-CNTL/PCI-OE/OE6/$1I296  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OE/OE6/$1I296/I0 ),
    .I1(NlwRenamedSig_OI_PCI_CMD10),
    .I2(\PCI-CNTL/LADX6 ),
    .I3(NlwRenamedSig_OI_CFG_HIT),
    .O(\PCI-CNTL/PCI-OE/OE6/NS_OE )
  );
  X_BUF   \PCI-CNTL/PCI-OE/OE5/$1I320  (
    .I(\PCI-CNTL/PCI-OE/OE5/Q ),
    .O(OE5)
  );
  X_BUF   \PCI-CNTL/PCI-OE/OE5/$1I311  (
    .I(\PCI-CNTL/END ),
    .O(\PCI-CNTL/PCI-OE/OE5/S )
  );
  X_BUF   \PCI-CNTL/PCI-OE/OE5/$1I310  (
    .I(\PCI-CNTL/PCI-OE/OE5/NS_OE ),
    .O(\PCI-CNTL/PCI-OE/OE5/R )
  );
  X_BUF   \PCI-CNTL/PCI-OE/OE5/$1I309  (
    .I(CLK),
    .O(\PCI-CNTL/PCI-OE/OE5/C )
  );
  X_AND2   \PCI-CNTL/PCI-OE/OE5/$1I307  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OE/OE5/$1I307/I0 ),
    .I1(\PCI-CNTL/PCI-OE/OE5/Q ),
    .O(\PCI-CNTL/PCI-OE/OE5/$1N301 )
  );
  X_OR2   \PCI-CNTL/PCI-OE/OE5/$1I306  (
    .I0(\PCI-CNTL/PCI-OE/OE5/S ),
    .I1(\PCI-CNTL/PCI-OE/OE5/$1N301 ),
    .O(\PCI-CNTL/PCI-OE/OE5/D )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-CNTL/PCI-OE/OE5/FDPE  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(\PCI-CNTL/PCI-OE/OE5/C ),
    .I(\PCI-CNTL/PCI-OE/OE5/D ),
    .O(\PCI-CNTL/PCI-OE/OE5/Q ),
    .RST(GND)
  );
  X_AND4   \PCI-CNTL/PCI-OE/OE5/$1I296  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OE/OE5/$1I296/I0 ),
    .I1(NlwRenamedSig_OI_PCI_CMD10),
    .I2(\PCI-CNTL/LADX5 ),
    .I3(NlwRenamedSig_OI_CFG_HIT),
    .O(\PCI-CNTL/PCI-OE/OE5/NS_OE )
  );
  X_BUF   \PCI-CNTL/PCI-OE/OE4/$1I320  (
    .I(\PCI-CNTL/PCI-OE/OE4/Q ),
    .O(OE4)
  );
  X_BUF   \PCI-CNTL/PCI-OE/OE4/$1I311  (
    .I(\PCI-CNTL/END ),
    .O(\PCI-CNTL/PCI-OE/OE4/S )
  );
  X_BUF   \PCI-CNTL/PCI-OE/OE4/$1I310  (
    .I(\PCI-CNTL/PCI-OE/OE4/NS_OE ),
    .O(\PCI-CNTL/PCI-OE/OE4/R )
  );
  X_BUF   \PCI-CNTL/PCI-OE/OE4/$1I309  (
    .I(CLK),
    .O(\PCI-CNTL/PCI-OE/OE4/C )
  );
  X_AND2   \PCI-CNTL/PCI-OE/OE4/$1I307  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OE/OE4/$1I307/I0 ),
    .I1(\PCI-CNTL/PCI-OE/OE4/Q ),
    .O(\PCI-CNTL/PCI-OE/OE4/$1N301 )
  );
  X_OR2   \PCI-CNTL/PCI-OE/OE4/$1I306  (
    .I0(\PCI-CNTL/PCI-OE/OE4/S ),
    .I1(\PCI-CNTL/PCI-OE/OE4/$1N301 ),
    .O(\PCI-CNTL/PCI-OE/OE4/D )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-CNTL/PCI-OE/OE4/FDPE  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(\PCI-CNTL/PCI-OE/OE4/C ),
    .I(\PCI-CNTL/PCI-OE/OE4/D ),
    .O(\PCI-CNTL/PCI-OE/OE4/Q ),
    .RST(GND)
  );
  X_AND4   \PCI-CNTL/PCI-OE/OE4/$1I296  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OE/OE4/$1I296/I0 ),
    .I1(NlwRenamedSig_OI_PCI_CMD10),
    .I2(\PCI-CNTL/LADX4 ),
    .I3(NlwRenamedSig_OI_CFG_HIT),
    .O(\PCI-CNTL/PCI-OE/OE4/NS_OE )
  );
  X_BUF   \PCI-CNTL/PCI-OE/OE3/$1I320  (
    .I(\PCI-CNTL/PCI-OE/OE3/Q ),
    .O(OE3)
  );
  X_BUF   \PCI-CNTL/PCI-OE/OE3/$1I311  (
    .I(\PCI-CNTL/END ),
    .O(\PCI-CNTL/PCI-OE/OE3/S )
  );
  X_BUF   \PCI-CNTL/PCI-OE/OE3/$1I310  (
    .I(\PCI-CNTL/PCI-OE/OE3/NS_OE ),
    .O(\PCI-CNTL/PCI-OE/OE3/R )
  );
  X_BUF   \PCI-CNTL/PCI-OE/OE3/$1I309  (
    .I(CLK),
    .O(\PCI-CNTL/PCI-OE/OE3/C )
  );
  X_AND2   \PCI-CNTL/PCI-OE/OE3/$1I307  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OE/OE3/$1I307/I0 ),
    .I1(\PCI-CNTL/PCI-OE/OE3/Q ),
    .O(\PCI-CNTL/PCI-OE/OE3/$1N301 )
  );
  X_OR2   \PCI-CNTL/PCI-OE/OE3/$1I306  (
    .I0(\PCI-CNTL/PCI-OE/OE3/S ),
    .I1(\PCI-CNTL/PCI-OE/OE3/$1N301 ),
    .O(\PCI-CNTL/PCI-OE/OE3/D )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-CNTL/PCI-OE/OE3/FDPE  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(\PCI-CNTL/PCI-OE/OE3/C ),
    .I(\PCI-CNTL/PCI-OE/OE3/D ),
    .O(\PCI-CNTL/PCI-OE/OE3/Q ),
    .RST(GND)
  );
  X_AND4   \PCI-CNTL/PCI-OE/OE3/$1I296  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OE/OE3/$1I296/I0 ),
    .I1(NlwRenamedSig_OI_PCI_CMD10),
    .I2(\PCI-CNTL/LADX3 ),
    .I3(NlwRenamedSig_OI_CFG_HIT),
    .O(\PCI-CNTL/PCI-OE/OE3/NS_OE )
  );
  X_BUF   \PCI-CNTL/PCI-OE/OE8/$1I320  (
    .I(\PCI-CNTL/PCI-OE/OE8/Q ),
    .O(OE8)
  );
  X_BUF   \PCI-CNTL/PCI-OE/OE8/$1I311  (
    .I(\PCI-CNTL/END ),
    .O(\PCI-CNTL/PCI-OE/OE8/S )
  );
  X_BUF   \PCI-CNTL/PCI-OE/OE8/$1I310  (
    .I(\PCI-CNTL/PCI-OE/OE8/NS_OE ),
    .O(\PCI-CNTL/PCI-OE/OE8/R )
  );
  X_BUF   \PCI-CNTL/PCI-OE/OE8/$1I309  (
    .I(CLK),
    .O(\PCI-CNTL/PCI-OE/OE8/C )
  );
  X_AND2   \PCI-CNTL/PCI-OE/OE8/$1I307  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OE/OE8/$1I307/I0 ),
    .I1(\PCI-CNTL/PCI-OE/OE8/Q ),
    .O(\PCI-CNTL/PCI-OE/OE8/$1N301 )
  );
  X_OR2   \PCI-CNTL/PCI-OE/OE8/$1I306  (
    .I0(\PCI-CNTL/PCI-OE/OE8/S ),
    .I1(\PCI-CNTL/PCI-OE/OE8/$1N301 ),
    .O(\PCI-CNTL/PCI-OE/OE8/D )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-CNTL/PCI-OE/OE8/FDPE  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(\PCI-CNTL/PCI-OE/OE8/C ),
    .I(\PCI-CNTL/PCI-OE/OE8/D ),
    .O(\PCI-CNTL/PCI-OE/OE8/Q ),
    .RST(GND)
  );
  X_AND4   \PCI-CNTL/PCI-OE/OE8/$1I296  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OE/OE8/$1I296/I0 ),
    .I1(NlwRenamedSig_OI_PCI_CMD10),
    .I2(\PCI-CNTL/LADX8 ),
    .I3(NlwRenamedSig_OI_CFG_HIT),
    .O(\PCI-CNTL/PCI-OE/OE8/NS_OE )
  );
  X_BUF   \PCI-CNTL/PCI-OE/OE9/$1I320  (
    .I(\PCI-CNTL/PCI-OE/OE9/Q ),
    .O(OE9)
  );
  X_BUF   \PCI-CNTL/PCI-OE/OE9/$1I311  (
    .I(\PCI-CNTL/END ),
    .O(\PCI-CNTL/PCI-OE/OE9/S )
  );
  X_BUF   \PCI-CNTL/PCI-OE/OE9/$1I310  (
    .I(\PCI-CNTL/PCI-OE/OE9/NS_OE ),
    .O(\PCI-CNTL/PCI-OE/OE9/R )
  );
  X_BUF   \PCI-CNTL/PCI-OE/OE9/$1I309  (
    .I(CLK),
    .O(\PCI-CNTL/PCI-OE/OE9/C )
  );
  X_AND2   \PCI-CNTL/PCI-OE/OE9/$1I307  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OE/OE9/$1I307/I0 ),
    .I1(\PCI-CNTL/PCI-OE/OE9/Q ),
    .O(\PCI-CNTL/PCI-OE/OE9/$1N301 )
  );
  X_OR2   \PCI-CNTL/PCI-OE/OE9/$1I306  (
    .I0(\PCI-CNTL/PCI-OE/OE9/S ),
    .I1(\PCI-CNTL/PCI-OE/OE9/$1N301 ),
    .O(\PCI-CNTL/PCI-OE/OE9/D )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-CNTL/PCI-OE/OE9/FDPE  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(\PCI-CNTL/PCI-OE/OE9/C ),
    .I(\PCI-CNTL/PCI-OE/OE9/D ),
    .O(\PCI-CNTL/PCI-OE/OE9/Q ),
    .RST(GND)
  );
  X_AND4   \PCI-CNTL/PCI-OE/OE9/$1I296  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OE/OE9/$1I296/I0 ),
    .I1(NlwRenamedSig_OI_PCI_CMD10),
    .I2(\PCI-CNTL/LADX9 ),
    .I3(NlwRenamedSig_OI_CFG_HIT),
    .O(\PCI-CNTL/PCI-OE/OE9/NS_OE )
  );
  X_BUF   \PCI-CNTL/PCI-OE/OE12/$1I320  (
    .I(\PCI-CNTL/PCI-OE/OE12/Q ),
    .O(OE12)
  );
  X_BUF   \PCI-CNTL/PCI-OE/OE12/$1I311  (
    .I(\PCI-CNTL/END ),
    .O(\PCI-CNTL/PCI-OE/OE12/S )
  );
  X_BUF   \PCI-CNTL/PCI-OE/OE12/$1I310  (
    .I(\PCI-CNTL/PCI-OE/OE12/NS_OE ),
    .O(\PCI-CNTL/PCI-OE/OE12/R )
  );
  X_BUF   \PCI-CNTL/PCI-OE/OE12/$1I309  (
    .I(CLK),
    .O(\PCI-CNTL/PCI-OE/OE12/C )
  );
  X_AND2   \PCI-CNTL/PCI-OE/OE12/$1I307  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OE/OE12/$1I307/I0 ),
    .I1(\PCI-CNTL/PCI-OE/OE12/Q ),
    .O(\PCI-CNTL/PCI-OE/OE12/$1N301 )
  );
  X_OR2   \PCI-CNTL/PCI-OE/OE12/$1I306  (
    .I0(\PCI-CNTL/PCI-OE/OE12/S ),
    .I1(\PCI-CNTL/PCI-OE/OE12/$1N301 ),
    .O(\PCI-CNTL/PCI-OE/OE12/D )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-CNTL/PCI-OE/OE12/FDPE  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(\PCI-CNTL/PCI-OE/OE12/C ),
    .I(\PCI-CNTL/PCI-OE/OE12/D ),
    .O(\PCI-CNTL/PCI-OE/OE12/Q ),
    .RST(GND)
  );
  X_AND4   \PCI-CNTL/PCI-OE/OE12/$1I296  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OE/OE12/$1I296/I0 ),
    .I1(NlwRenamedSig_OI_PCI_CMD10),
    .I2(\PCI-CNTL/LADX12 ),
    .I3(NlwRenamedSig_OI_CFG_HIT),
    .O(\PCI-CNTL/PCI-OE/OE12/NS_OE )
  );
  X_BUF   \PCI-CNTL/PCI-OE/OE1/$1I320  (
    .I(\PCI-CNTL/PCI-OE/OE1/Q ),
    .O(OE1)
  );
  X_BUF   \PCI-CNTL/PCI-OE/OE1/$1I311  (
    .I(\PCI-CNTL/END ),
    .O(\PCI-CNTL/PCI-OE/OE1/S )
  );
  X_BUF   \PCI-CNTL/PCI-OE/OE1/$1I310  (
    .I(\PCI-CNTL/PCI-OE/OE1/NS_OE ),
    .O(\PCI-CNTL/PCI-OE/OE1/R )
  );
  X_BUF   \PCI-CNTL/PCI-OE/OE1/$1I309  (
    .I(CLK),
    .O(\PCI-CNTL/PCI-OE/OE1/C )
  );
  X_AND2   \PCI-CNTL/PCI-OE/OE1/$1I307  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OE/OE1/$1I307/I0 ),
    .I1(\PCI-CNTL/PCI-OE/OE1/Q ),
    .O(\PCI-CNTL/PCI-OE/OE1/$1N301 )
  );
  X_OR2   \PCI-CNTL/PCI-OE/OE1/$1I306  (
    .I0(\PCI-CNTL/PCI-OE/OE1/S ),
    .I1(\PCI-CNTL/PCI-OE/OE1/$1N301 ),
    .O(\PCI-CNTL/PCI-OE/OE1/D )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-CNTL/PCI-OE/OE1/FDPE  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(\PCI-CNTL/PCI-OE/OE1/C ),
    .I(\PCI-CNTL/PCI-OE/OE1/D ),
    .O(\PCI-CNTL/PCI-OE/OE1/Q ),
    .RST(GND)
  );
  X_AND4   \PCI-CNTL/PCI-OE/OE1/$1I296  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OE/OE1/$1I296/I0 ),
    .I1(NlwRenamedSig_OI_PCI_CMD10),
    .I2(\PCI-CNTL/LADX1 ),
    .I3(NlwRenamedSig_OI_CFG_HIT),
    .O(\PCI-CNTL/PCI-OE/OE1/NS_OE )
  );
  X_ZERO   \PCI-CNTL/PCI-OE/$1I849/$1I2218  (
    .O(\PCI-CNTL/PCI-OE/$1I849/$1N2216 )
  );
  X_BUF   \PCI-CNTL/PCI-OE/$1I849/NS  (
    .I(\PCI-CNTL/PCI-OE/$1I849/$1N2216 ),
    .O(OE13)
  );
  X_ZERO   \PCI-CNTL/PCI-OE/$1I850/$1I2218  (
    .O(\PCI-CNTL/PCI-OE/$1I850/$1N2216 )
  );
  X_BUF   \PCI-CNTL/PCI-OE/$1I850/NS  (
    .I(\PCI-CNTL/PCI-OE/$1I850/$1N2216 ),
    .O(OE0)
  );
  X_ZERO   \PCI-CNTL/PCI-OE/$1I853/$1I2218  (
    .O(\PCI-CNTL/PCI-OE/$1I853/$1N2216 )
  );
  X_BUF   \PCI-CNTL/PCI-OE/$1I853/NS  (
    .I(\PCI-CNTL/PCI-OE/$1I853/$1N2216 ),
    .O(OE2)
  );
  X_ZERO   \PCI-CNTL/PCI-OE/$1I868/$1I2218  (
    .O(\PCI-CNTL/PCI-OE/$1I868/$1N2216 )
  );
  X_BUF   \PCI-CNTL/PCI-OE/$1I868/NS  (
    .I(\PCI-CNTL/PCI-OE/$1I868/$1N2216 ),
    .O(OE11)
  );
  X_ZERO   \PCI-CNTL/PCI-OE/$1I870/$1I2218  (
    .O(\PCI-CNTL/PCI-OE/$1I870/$1N2216 )
  );
  X_BUF   \PCI-CNTL/PCI-OE/$1I870/NS  (
    .I(\PCI-CNTL/PCI-OE/$1I870/$1N2216 ),
    .O(OE14)
  );
  X_ZERO   \PCI-CNTL/PCI-OE/$1I872/$1I2218  (
    .O(\PCI-CNTL/PCI-OE/$1I872/$1N2216 )
  );
  X_BUF   \PCI-CNTL/PCI-OE/$1I872/NS  (
    .I(\PCI-CNTL/PCI-OE/$1I872/$1N2216 ),
    .O(OE10)
  );
  X_AND4   \PCI-CNTL/PCI-OE/DEC-F/AND4  (
    .I0(NlwRenamedSig_OI_ADDR2),
    .I1(NlwRenamedSig_OI_ADDR3),
    .I2(NlwRenamedSig_OI_ADDR4),
    .I3(NlwRenamedSig_OI_ADDR5),
    .O(\PCI-CNTL/PCI-OE/3CH )
  );
  X_AND4   \PCI-CNTL/PCI-OE/DEC-E/AND4  (
    .I0(\PCI-CNTL/PCI-OE/DEC-E/$1N2275 ),
    .I1(NlwRenamedSig_OI_ADDR3),
    .I2(NlwRenamedSig_OI_ADDR4),
    .I3(NlwRenamedSig_OI_ADDR5),
    .O(\PCI-CNTL/PCI-OE/38H )
  );
  X_INV   \PCI-CNTL/PCI-OE/DEC-E/INV0  (
    .I(NlwRenamedSig_OI_ADDR2),
    .O(\PCI-CNTL/PCI-OE/DEC-E/$1N2275 )
  );
  X_AND4   \PCI-CNTL/PCI-OE/DEC-D/AND4  (
    .I0(NlwRenamedSig_OI_ADDR2),
    .I1(\PCI-CNTL/PCI-OE/DEC-D/$1N2290 ),
    .I2(NlwRenamedSig_OI_ADDR4),
    .I3(NlwRenamedSig_OI_ADDR5),
    .O(\PCI-CNTL/PCI-OE/34H )
  );
  X_INV   \PCI-CNTL/PCI-OE/DEC-D/INV1  (
    .I(NlwRenamedSig_OI_ADDR3),
    .O(\PCI-CNTL/PCI-OE/DEC-D/$1N2290 )
  );
  X_AND4   \PCI-CNTL/PCI-OE/DEC-C/AND4  (
    .I0(\PCI-CNTL/PCI-OE/DEC-C/$1N2289 ),
    .I1(\PCI-CNTL/PCI-OE/DEC-C/$1N2290 ),
    .I2(NlwRenamedSig_OI_ADDR4),
    .I3(NlwRenamedSig_OI_ADDR5),
    .O(\PCI-CNTL/PCI-OE/30H )
  );
  X_INV   \PCI-CNTL/PCI-OE/DEC-C/INV1  (
    .I(NlwRenamedSig_OI_ADDR3),
    .O(\PCI-CNTL/PCI-OE/DEC-C/$1N2290 )
  );
  X_INV   \PCI-CNTL/PCI-OE/DEC-C/INV0  (
    .I(NlwRenamedSig_OI_ADDR2),
    .O(\PCI-CNTL/PCI-OE/DEC-C/$1N2289 )
  );
  X_AND4   \PCI-CNTL/PCI-OE/DEC-9/AND4  (
    .I0(NlwRenamedSig_OI_ADDR2),
    .I1(\PCI-CNTL/PCI-OE/DEC-9/$1N2276 ),
    .I2(\PCI-CNTL/PCI-OE/DEC-9/$1N2277 ),
    .I3(NlwRenamedSig_OI_ADDR5),
    .O(\PCI-CNTL/PCI-OE/24H )
  );
  X_INV   \PCI-CNTL/PCI-OE/DEC-9/INV2  (
    .I(NlwRenamedSig_OI_ADDR4),
    .O(\PCI-CNTL/PCI-OE/DEC-9/$1N2277 )
  );
  X_INV   \PCI-CNTL/PCI-OE/DEC-9/INV1  (
    .I(NlwRenamedSig_OI_ADDR3),
    .O(\PCI-CNTL/PCI-OE/DEC-9/$1N2276 )
  );
  X_AND4   \PCI-CNTL/PCI-OE/DEC-8/AND4  (
    .I0(\PCI-CNTL/PCI-OE/DEC-8/$1N2275 ),
    .I1(\PCI-CNTL/PCI-OE/DEC-8/$1N2276 ),
    .I2(\PCI-CNTL/PCI-OE/DEC-8/$1N2277 ),
    .I3(NlwRenamedSig_OI_ADDR5),
    .O(\PCI-CNTL/PCI-OE/20H )
  );
  X_INV   \PCI-CNTL/PCI-OE/DEC-8/INV2  (
    .I(NlwRenamedSig_OI_ADDR4),
    .O(\PCI-CNTL/PCI-OE/DEC-8/$1N2277 )
  );
  X_INV   \PCI-CNTL/PCI-OE/DEC-8/INV1  (
    .I(NlwRenamedSig_OI_ADDR3),
    .O(\PCI-CNTL/PCI-OE/DEC-8/$1N2276 )
  );
  X_INV   \PCI-CNTL/PCI-OE/DEC-8/INV0  (
    .I(NlwRenamedSig_OI_ADDR2),
    .O(\PCI-CNTL/PCI-OE/DEC-8/$1N2275 )
  );
  X_AND4   \PCI-CNTL/PCI-OE/DEC-7/AND4  (
    .I0(NlwRenamedSig_OI_ADDR2),
    .I1(NlwRenamedSig_OI_ADDR3),
    .I2(NlwRenamedSig_OI_ADDR4),
    .I3(\PCI-CNTL/PCI-OE/DEC-7/$1N2283 ),
    .O(\PCI-CNTL/PCI-OE/1CH )
  );
  X_INV   \PCI-CNTL/PCI-OE/DEC-7/INV3  (
    .I(NlwRenamedSig_OI_ADDR5),
    .O(\PCI-CNTL/PCI-OE/DEC-7/$1N2283 )
  );
  X_AND4   \PCI-CNTL/PCI-OE/DEC-6/AND4  (
    .I0(\PCI-CNTL/PCI-OE/DEC-6/$1N2275 ),
    .I1(NlwRenamedSig_OI_ADDR3),
    .I2(NlwRenamedSig_OI_ADDR4),
    .I3(\PCI-CNTL/PCI-OE/DEC-6/$1N2283 ),
    .O(\PCI-CNTL/PCI-OE/18H )
  );
  X_INV   \PCI-CNTL/PCI-OE/DEC-6/INV3  (
    .I(NlwRenamedSig_OI_ADDR5),
    .O(\PCI-CNTL/PCI-OE/DEC-6/$1N2283 )
  );
  X_INV   \PCI-CNTL/PCI-OE/DEC-6/INV0  (
    .I(NlwRenamedSig_OI_ADDR2),
    .O(\PCI-CNTL/PCI-OE/DEC-6/$1N2275 )
  );
  X_AND4   \PCI-CNTL/PCI-OE/DEC-B/AND4  (
    .I0(NlwRenamedSig_OI_ADDR2),
    .I1(NlwRenamedSig_OI_ADDR3),
    .I2(\PCI-CNTL/PCI-OE/DEC-B/$1N2277 ),
    .I3(NlwRenamedSig_OI_ADDR5),
    .O(\PCI-CNTL/PCI-OE/2CH )
  );
  X_INV   \PCI-CNTL/PCI-OE/DEC-B/INV2  (
    .I(NlwRenamedSig_OI_ADDR4),
    .O(\PCI-CNTL/PCI-OE/DEC-B/$1N2277 )
  );
  X_AND4   \PCI-CNTL/PCI-OE/DEC-A/AND4  (
    .I0(\PCI-CNTL/PCI-OE/DEC-A/$1N2275 ),
    .I1(NlwRenamedSig_OI_ADDR3),
    .I2(\PCI-CNTL/PCI-OE/DEC-A/$1N2277 ),
    .I3(NlwRenamedSig_OI_ADDR5),
    .O(\PCI-CNTL/PCI-OE/28H )
  );
  X_INV   \PCI-CNTL/PCI-OE/DEC-A/INV2  (
    .I(NlwRenamedSig_OI_ADDR4),
    .O(\PCI-CNTL/PCI-OE/DEC-A/$1N2277 )
  );
  X_INV   \PCI-CNTL/PCI-OE/DEC-A/INV0  (
    .I(NlwRenamedSig_OI_ADDR2),
    .O(\PCI-CNTL/PCI-OE/DEC-A/$1N2275 )
  );
  X_AND4   \PCI-CNTL/PCI-OE/DEC-3/AND4  (
    .I0(NlwRenamedSig_OI_ADDR2),
    .I1(NlwRenamedSig_OI_ADDR3),
    .I2(\PCI-CNTL/PCI-OE/DEC-3/$1N2277 ),
    .I3(\PCI-CNTL/PCI-OE/DEC-3/$1N2283 ),
    .O(\PCI-CNTL/PCI-OE/0CH )
  );
  X_INV   \PCI-CNTL/PCI-OE/DEC-3/INV3  (
    .I(NlwRenamedSig_OI_ADDR5),
    .O(\PCI-CNTL/PCI-OE/DEC-3/$1N2283 )
  );
  X_INV   \PCI-CNTL/PCI-OE/DEC-3/INV2  (
    .I(NlwRenamedSig_OI_ADDR4),
    .O(\PCI-CNTL/PCI-OE/DEC-3/$1N2277 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-CNTL/PCI-OE/$2I617/FDPE  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(CLK),
    .I(\PCI-CNTL/PCI-OE/$2I617/D ),
    .O(OE_ROM),
    .RST(GND)
  );
  X_OR2   \PCI-CNTL/PCI-OE/$2I617/$1I12  (
    .I0(\PCI-CNTL/END ),
    .I1(\PCI-CNTL/PCI-OE/$2I617/$1N18 ),
    .O(\PCI-CNTL/PCI-OE/$2I617/D )
  );
  X_AND2   \PCI-CNTL/PCI-OE/$2I617/$1I11  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OE/$2I617/$1I11/I0 ),
    .I1(OE_ROM),
    .O(\PCI-CNTL/PCI-OE/$2I617/$1N18 )
  );
  X_OR4   \PCI-CNTL/PCI-OE/OR16/G3  (
    .I0(\PCI-CNTL/PCI-OE/$2N747 ),
    .I1(\PCI-CNTL/PCI-OE/$2N746 ),
    .I2(\PCI-CNTL/PCI-OE/$2N745 ),
    .I3(\PCI-CNTL/PCI-OE/$2N744 ),
    .O(\PCI-CNTL/PCI-OE/OR16/$1N2234 )
  );
  X_OR4   \PCI-CNTL/PCI-OE/OR16/G2  (
    .I0(\PCI-CNTL/PCI-OE/$2N751 ),
    .I1(\PCI-CNTL/PCI-OE/$2N750 ),
    .I2(\PCI-CNTL/PCI-OE/$2N749 ),
    .I3(\PCI-CNTL/PCI-OE/$2N748 ),
    .O(\PCI-CNTL/PCI-OE/OR16/$1N2243 )
  );
  X_OR4   \PCI-CNTL/PCI-OE/OR16/O  (
    .I0(\PCI-CNTL/PCI-OE/OR16/$1N2216 ),
    .I1(\PCI-CNTL/PCI-OE/OR16/$1N2224 ),
    .I2(\PCI-CNTL/PCI-OE/OR16/$1N2243 ),
    .I3(\PCI-CNTL/PCI-OE/OR16/$1N2234 ),
    .O(\PCI-CNTL/PCI-OE/X )
  );
  X_OR4   \PCI-CNTL/PCI-OE/OR16/G1  (
    .I0(\PCI-CNTL/PCI-OE/$2N755 ),
    .I1(\PCI-CNTL/PCI-OE/$2N754 ),
    .I2(\PCI-CNTL/PCI-OE/$2N753 ),
    .I3(\PCI-CNTL/PCI-OE/$2N752 ),
    .O(\PCI-CNTL/PCI-OE/OR16/$1N2224 )
  );
  X_OR4   \PCI-CNTL/PCI-OE/OR16/G0  (
    .I0(\PCI-CNTL/PCI-OE/$2N697 ),
    .I1(\PCI-CNTL/PCI-OE/$2N758 ),
    .I2(\PCI-CNTL/PCI-OE/$2N757 ),
    .I3(\PCI-CNTL/PCI-OE/$2N756 ),
    .O(\PCI-CNTL/PCI-OE/OR16/$1N2216 )
  );
  X_AND4   \PCI-CNTL/PCI-OE/DEC-5/AND4  (
    .I0(NlwRenamedSig_OI_ADDR2),
    .I1(\PCI-CNTL/PCI-OE/DEC-5/$1N2276 ),
    .I2(NlwRenamedSig_OI_ADDR4),
    .I3(\PCI-CNTL/PCI-OE/DEC-5/$1N2283 ),
    .O(\PCI-CNTL/PCI-OE/14H )
  );
  X_INV   \PCI-CNTL/PCI-OE/DEC-5/INV3  (
    .I(NlwRenamedSig_OI_ADDR5),
    .O(\PCI-CNTL/PCI-OE/DEC-5/$1N2283 )
  );
  X_INV   \PCI-CNTL/PCI-OE/DEC-5/INV1  (
    .I(NlwRenamedSig_OI_ADDR3),
    .O(\PCI-CNTL/PCI-OE/DEC-5/$1N2276 )
  );
  X_AND4   \PCI-CNTL/PCI-OE/DEC-4/AND4  (
    .I0(\PCI-CNTL/PCI-OE/DEC-4/$1N2275 ),
    .I1(\PCI-CNTL/PCI-OE/DEC-4/$1N2276 ),
    .I2(NlwRenamedSig_OI_ADDR4),
    .I3(\PCI-CNTL/PCI-OE/DEC-4/$1N2283 ),
    .O(\PCI-CNTL/PCI-OE/10H )
  );
  X_INV   \PCI-CNTL/PCI-OE/DEC-4/INV3  (
    .I(NlwRenamedSig_OI_ADDR5),
    .O(\PCI-CNTL/PCI-OE/DEC-4/$1N2283 )
  );
  X_INV   \PCI-CNTL/PCI-OE/DEC-4/INV1  (
    .I(NlwRenamedSig_OI_ADDR3),
    .O(\PCI-CNTL/PCI-OE/DEC-4/$1N2276 )
  );
  X_INV   \PCI-CNTL/PCI-OE/DEC-4/INV0  (
    .I(NlwRenamedSig_OI_ADDR2),
    .O(\PCI-CNTL/PCI-OE/DEC-4/$1N2275 )
  );
  X_AND4   \PCI-CNTL/PCI-OE/DEC-2/AND4  (
    .I0(\PCI-CNTL/PCI-OE/DEC-2/$1N2275 ),
    .I1(NlwRenamedSig_OI_ADDR3),
    .I2(\PCI-CNTL/PCI-OE/DEC-2/$1N2277 ),
    .I3(\PCI-CNTL/PCI-OE/DEC-2/$1N2283 ),
    .O(\PCI-CNTL/PCI-OE/08H )
  );
  X_INV   \PCI-CNTL/PCI-OE/DEC-2/INV3  (
    .I(NlwRenamedSig_OI_ADDR5),
    .O(\PCI-CNTL/PCI-OE/DEC-2/$1N2283 )
  );
  X_INV   \PCI-CNTL/PCI-OE/DEC-2/INV2  (
    .I(NlwRenamedSig_OI_ADDR4),
    .O(\PCI-CNTL/PCI-OE/DEC-2/$1N2277 )
  );
  X_INV   \PCI-CNTL/PCI-OE/DEC-2/INV0  (
    .I(NlwRenamedSig_OI_ADDR2),
    .O(\PCI-CNTL/PCI-OE/DEC-2/$1N2275 )
  );
  X_INV   \PCI-CNTL/PCI-OE/DEC-1/INV1  (
    .I(NlwRenamedSig_OI_ADDR3),
    .O(\PCI-CNTL/PCI-OE/DEC-1/$1N2280 )
  );
  X_INV   \PCI-CNTL/PCI-OE/DEC-1/INV2  (
    .I(NlwRenamedSig_OI_ADDR4),
    .O(\PCI-CNTL/PCI-OE/DEC-1/$1N2278 )
  );
  X_INV   \PCI-CNTL/PCI-OE/DEC-1/INV3  (
    .I(NlwRenamedSig_OI_ADDR5),
    .O(\PCI-CNTL/PCI-OE/DEC-1/$1N2277 )
  );
  X_AND4   \PCI-CNTL/PCI-OE/DEC-1/AND4  (
    .I0(NlwRenamedSig_OI_ADDR2),
    .I1(\PCI-CNTL/PCI-OE/DEC-1/$1N2280 ),
    .I2(\PCI-CNTL/PCI-OE/DEC-1/$1N2278 ),
    .I3(\PCI-CNTL/PCI-OE/DEC-1/$1N2277 ),
    .O(\PCI-CNTL/PCI-OE/04H )
  );
  X_AND4   \PCI-CNTL/PCI-OE/DEC-0/AND4  (
    .I0(\PCI-CNTL/PCI-OE/DEC-0/$1N2275 ),
    .I1(\PCI-CNTL/PCI-OE/DEC-0/$1N2276 ),
    .I2(\PCI-CNTL/PCI-OE/DEC-0/$1N2277 ),
    .I3(\PCI-CNTL/PCI-OE/DEC-0/$1N2283 ),
    .O(\PCI-CNTL/PCI-OE/00H )
  );
  X_INV   \PCI-CNTL/PCI-OE/DEC-0/INV3  (
    .I(NlwRenamedSig_OI_ADDR5),
    .O(\PCI-CNTL/PCI-OE/DEC-0/$1N2283 )
  );
  X_INV   \PCI-CNTL/PCI-OE/DEC-0/INV2  (
    .I(NlwRenamedSig_OI_ADDR4),
    .O(\PCI-CNTL/PCI-OE/DEC-0/$1N2277 )
  );
  X_INV   \PCI-CNTL/PCI-OE/DEC-0/INV1  (
    .I(NlwRenamedSig_OI_ADDR3),
    .O(\PCI-CNTL/PCI-OE/DEC-0/$1N2276 )
  );
  X_INV   \PCI-CNTL/PCI-OE/DEC-0/INV0  (
    .I(NlwRenamedSig_OI_ADDR2),
    .O(\PCI-CNTL/PCI-OE/DEC-0/$1N2275 )
  );
  X_BUF   \PCI-CNTL/PCI-OE/SW1/$1I2289/NC  (
    .I(\PCI-CNTL/PCI-OE/04H ),
    .O(\NLW_PCI-CNTL/PCI-OE/SW1/$1I2289/NC_O_UNCONNECTED )
  );
  X_ZERO   \PCI-CNTL/PCI-OE/SW1/$1I2290/$1I2218  (
    .O(\PCI-CNTL/PCI-OE/SW1/$1I2290/$1N2216 )
  );
  X_BUF   \PCI-CNTL/PCI-OE/SW1/$1I2290/NS  (
    .I(\PCI-CNTL/PCI-OE/SW1/$1I2290/$1N2216 ),
    .O(\PCI-CNTL/PCI-OE/$2N758 )
  );
  X_BUF   \PCI-CNTL/PCI-OE/SW7/$1I2293  (
    .I(\PCI-CNTL/PCI-OE/1CH ),
    .O(\PCI-CNTL/PCI-OE/$2N752 )
  );
  X_BUF   \PCI-CNTL/PCI-OE/SW8/$1I2293  (
    .I(\PCI-CNTL/PCI-OE/20H ),
    .O(\PCI-CNTL/PCI-OE/$2N751 )
  );
  X_BUF   \PCI-CNTL/PCI-OE/SW9/$1I2293  (
    .I(\PCI-CNTL/PCI-OE/24H ),
    .O(\PCI-CNTL/PCI-OE/$2N750 )
  );
  X_BUF   \PCI-CNTL/PCI-OE/SW10/$1I2293  (
    .I(\PCI-CNTL/PCI-OE/28H ),
    .O(\PCI-CNTL/PCI-OE/$2N749 )
  );
  X_BUF   \PCI-CNTL/PCI-OE/SW12/$1I2293  (
    .I(\PCI-CNTL/PCI-OE/30H ),
    .O(\PCI-CNTL/PCI-OE/$2N747 )
  );
  X_BUF   \PCI-CNTL/PCI-OE/SW14/$1I2293  (
    .I(\PCI-CNTL/PCI-OE/38H ),
    .O(\PCI-CNTL/PCI-OE/$2N745 )
  );
  X_BUF   \PCI-CNTL/PCI-OE/SW15/$1I2289/NC  (
    .I(\PCI-CNTL/PCI-OE/3CH ),
    .O(\NLW_PCI-CNTL/PCI-OE/SW15/$1I2289/NC_O_UNCONNECTED )
  );
  X_ZERO   \PCI-CNTL/PCI-OE/SW15/$1I2290/$1I2218  (
    .O(\PCI-CNTL/PCI-OE/SW15/$1I2290/$1N2216 )
  );
  X_BUF   \PCI-CNTL/PCI-OE/SW15/$1I2290/NS  (
    .I(\PCI-CNTL/PCI-OE/SW15/$1I2290/$1N2216 ),
    .O(\PCI-CNTL/PCI-OE/$2N744 )
  );
  X_BUF   \PCI-CNTL/PCI-OE/SW0/$1I2293  (
    .I(\PCI-CNTL/PCI-OE/00H ),
    .O(\PCI-CNTL/PCI-OE/$2N697 )
  );
  X_BUF   \PCI-CNTL/PCI-OE/SW2/$1I2293  (
    .I(\PCI-CNTL/PCI-OE/08H ),
    .O(\PCI-CNTL/PCI-OE/$2N757 )
  );
  X_BUF   \PCI-CNTL/PCI-OE/SW3/$1I2289/NC  (
    .I(\PCI-CNTL/PCI-OE/0CH ),
    .O(\NLW_PCI-CNTL/PCI-OE/SW3/$1I2289/NC_O_UNCONNECTED )
  );
  X_ZERO   \PCI-CNTL/PCI-OE/SW3/$1I2290/$1I2218  (
    .O(\PCI-CNTL/PCI-OE/SW3/$1I2290/$1N2216 )
  );
  X_BUF   \PCI-CNTL/PCI-OE/SW3/$1I2290/NS  (
    .I(\PCI-CNTL/PCI-OE/SW3/$1I2290/$1N2216 ),
    .O(\PCI-CNTL/PCI-OE/$2N756 )
  );
  X_BUF   \PCI-CNTL/PCI-OE/SW11/$1I2293  (
    .I(\PCI-CNTL/PCI-OE/2CH ),
    .O(\PCI-CNTL/PCI-OE/$2N748 )
  );
  X_BUF   \PCI-CNTL/PCI-OE/SW13/$1I2293  (
    .I(\PCI-CNTL/PCI-OE/34H ),
    .O(\PCI-CNTL/PCI-OE/$2N746 )
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE15/G0  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N0 ),
    .I3(\PCI-CNTL/LADX15 ),
    .O(CE15_0)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE15/G1  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N1 ),
    .I3(\PCI-CNTL/LADX15 ),
    .O(CE15_1)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE15/G2  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N2 ),
    .I3(\PCI-CNTL/LADX15 ),
    .O(CE15_2)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE15/G3  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N3 ),
    .I3(\PCI-CNTL/LADX15 ),
    .O(CE15_3)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE14/G0  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N0 ),
    .I3(\PCI-CNTL/LADX14 ),
    .O(CE14_0)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE14/G1  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N1 ),
    .I3(\PCI-CNTL/LADX14 ),
    .O(CE14_1)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE14/G2  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N2 ),
    .I3(\PCI-CNTL/LADX14 ),
    .O(CE14_2)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE14/G3  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N3 ),
    .I3(\PCI-CNTL/LADX14 ),
    .O(CE14_3)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE13/G0  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N0 ),
    .I3(\PCI-CNTL/LADX13 ),
    .O(CE13_0)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE13/G1  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N1 ),
    .I3(\PCI-CNTL/LADX13 ),
    .O(CE13_1)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE13/G2  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N2 ),
    .I3(\PCI-CNTL/LADX13 ),
    .O(CE13_2)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE13/G3  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N3 ),
    .I3(\PCI-CNTL/LADX13 ),
    .O(CE13_3)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE12/G0  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N0 ),
    .I3(\PCI-CNTL/LADX12 ),
    .O(CE12_0)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE12/G1  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N1 ),
    .I3(\PCI-CNTL/LADX12 ),
    .O(CE12_1)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE12/G2  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N2 ),
    .I3(\PCI-CNTL/LADX12 ),
    .O(CE12_2)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE12/G3  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N3 ),
    .I3(\PCI-CNTL/LADX12 ),
    .O(CE12_3)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE8/G0  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N0 ),
    .I3(\PCI-CNTL/LADX8 ),
    .O(CE8_0)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE8/G1  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N1 ),
    .I3(\PCI-CNTL/LADX8 ),
    .O(CE8_1)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE8/G2  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N2 ),
    .I3(\PCI-CNTL/LADX8 ),
    .O(CE8_2)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE8/G3  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N3 ),
    .I3(\PCI-CNTL/LADX8 ),
    .O(CE8_3)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE9/G0  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N0 ),
    .I3(\PCI-CNTL/LADX9 ),
    .O(CE9_0)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE9/G1  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N1 ),
    .I3(\PCI-CNTL/LADX9 ),
    .O(CE9_1)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE9/G2  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N2 ),
    .I3(\PCI-CNTL/LADX9 ),
    .O(CE9_2)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE9/G3  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N3 ),
    .I3(\PCI-CNTL/LADX9 ),
    .O(CE9_3)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE10/G0  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N0 ),
    .I3(\PCI-CNTL/LADX10 ),
    .O(CE10_0)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE10/G1  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N1 ),
    .I3(\PCI-CNTL/LADX10 ),
    .O(CE10_1)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE10/G2  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N2 ),
    .I3(\PCI-CNTL/LADX10 ),
    .O(CE10_2)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE10/G3  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N3 ),
    .I3(\PCI-CNTL/LADX10 ),
    .O(CE10_3)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE11/G0  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N0 ),
    .I3(\PCI-CNTL/LADX11 ),
    .O(CE11_0)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE11/G1  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N1 ),
    .I3(\PCI-CNTL/LADX11 ),
    .O(CE11_1)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE11/G2  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N2 ),
    .I3(\PCI-CNTL/LADX11 ),
    .O(CE11_2)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE11/G3  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N3 ),
    .I3(\PCI-CNTL/LADX11 ),
    .O(CE11_3)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE4/G0  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N0 ),
    .I3(\PCI-CNTL/LADX4 ),
    .O(CE4_0)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE4/G1  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N1 ),
    .I3(\PCI-CNTL/LADX4 ),
    .O(CE4_1)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE4/G2  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N2 ),
    .I3(\PCI-CNTL/LADX4 ),
    .O(CE4_2)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE4/G3  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N3 ),
    .I3(\PCI-CNTL/LADX4 ),
    .O(CE4_3)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE5/G0  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N0 ),
    .I3(\PCI-CNTL/LADX5 ),
    .O(CE5_0)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE5/G1  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N1 ),
    .I3(\PCI-CNTL/LADX5 ),
    .O(CE5_1)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE5/G2  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N2 ),
    .I3(\PCI-CNTL/LADX5 ),
    .O(CE5_2)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE5/G3  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N3 ),
    .I3(\PCI-CNTL/LADX5 ),
    .O(CE5_3)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE6/G0  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N0 ),
    .I3(\PCI-CNTL/LADX6 ),
    .O(CE6_0)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE6/G1  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N1 ),
    .I3(\PCI-CNTL/LADX6 ),
    .O(CE6_1)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE6/G2  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N2 ),
    .I3(\PCI-CNTL/LADX6 ),
    .O(CE6_2)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE6/G3  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N3 ),
    .I3(\PCI-CNTL/LADX6 ),
    .O(CE6_3)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE7/G0  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N0 ),
    .I3(\PCI-CNTL/LADX7 ),
    .O(CE7_0)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE7/G1  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N1 ),
    .I3(\PCI-CNTL/LADX7 ),
    .O(CE7_1)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE7/G2  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N2 ),
    .I3(\PCI-CNTL/LADX7 ),
    .O(CE7_2)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE7/G3  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N3 ),
    .I3(\PCI-CNTL/LADX7 ),
    .O(CE7_3)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE0/G0  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N0 ),
    .I3(\PCI-CNTL/LADX0 ),
    .O(CE0_0)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE0/G1  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N1 ),
    .I3(\PCI-CNTL/LADX0 ),
    .O(CE0_1)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE0/G2  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N2 ),
    .I3(\PCI-CNTL/LADX0 ),
    .O(CE0_2)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE0/G3  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N3 ),
    .I3(\PCI-CNTL/LADX0 ),
    .O(CE0_3)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE1/G0  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N0 ),
    .I3(\PCI-CNTL/LADX1 ),
    .O(CE1_0)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE1/G1  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N1 ),
    .I3(\PCI-CNTL/LADX1 ),
    .O(CE1_1)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE1/G2  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N2 ),
    .I3(\PCI-CNTL/LADX1 ),
    .O(CE1_2)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE1/G3  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N3 ),
    .I3(\PCI-CNTL/LADX1 ),
    .O(CE1_3)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE2/G0  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N0 ),
    .I3(\PCI-CNTL/LADX2 ),
    .O(CE2_0)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE2/G1  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N1 ),
    .I3(\PCI-CNTL/LADX2 ),
    .O(CE2_1)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE2/G2  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N2 ),
    .I3(\PCI-CNTL/LADX2 ),
    .O(CE2_2)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE2/G3  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N3 ),
    .I3(\PCI-CNTL/LADX2 ),
    .O(CE2_3)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE3/G0  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N0 ),
    .I3(\PCI-CNTL/LADX3 ),
    .O(CE3_0)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE3/G1  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N1 ),
    .I3(\PCI-CNTL/LADX3 ),
    .O(CE3_1)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE3/G2  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N2 ),
    .I3(\PCI-CNTL/LADX3 ),
    .O(CE3_2)
  );
  X_AND4   \PCI-CNTL/PCI-CE/CE3/G3  (
    .I0(\PCI-CNTL/DSTR ),
    .I1(NlwRenamedSig_OI_PCI_CMD11),
    .I2(\PCI-CNTL/CBE_N3 ),
    .I3(\PCI-CNTL/LADX3 ),
    .O(CE3_3)
  );
  X_BUF   \PCI-CNTL/$1I972/NC  (
    .I(SLOT64),
    .O(\NLW_PCI-CNTL/$1I972/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-CNTL/$1I974/NC  (
    .I(CFG115),
    .O(\NLW_PCI-CNTL/$1I974/NC_O_UNCONNECTED )
  );
  X_OR2   \PCI-CNTL/$1I995/$1I2214  (
    .I0(\PCI-CNTL/$1N1000 ),
    .I1(\PCI-CNTL/HOLD_APERR ),
    .O(\PCI-CNTL/$1I995/$1N2215 )
  );
  X_AND2   \PCI-CNTL/$1I995/$1I2213  (
    .I0(\NlwInverterSignal_PCI-CNTL/$1I995/$1I2213/I0 ),
    .I1(\PCI-CNTL/$1I995/$1N2215 ),
    .O(\PCI-CNTL/$1I995/D )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/$1I995/FDCE  (
    .CE(VCC),
    .CLK(CLK),
    .I(\PCI-CNTL/$1I995/D ),
    .O(\PCI-CNTL/HOLD_APERR ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-CNTL/PCI-TSM/PCI-IDLE/IDLE1_FF  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(CLK),
    .I(\PCI-CNTL/PCI-TSM/PCI-IDLE/NS_IDLE ),
    .O(IDLE_DUP),
    .RST(GND)
  );
  X_AND2   \PCI-CNTL/PCI-TSM/PCI-IDLE/$1I498  (
    .I0(\FRAME- ),
    .I1(BACKOFF_INT),
    .O(\PCI-CNTL/PCI-TSM/PCI-IDLE/BKOF_NS_TNAR )
  );
  X_OR2   \PCI-CNTL/PCI-TSM/PCI-IDLE/$1I497  (
    .I0(\PCI-CNTL/PCI-TSM/PCI-IDLE/BKOF_NS_TNAR ),
    .I1(\PCI-CNTL/PCI-TSM/PCI-IDLE/DATA_NS_TNAR ),
    .O(\PCI-CNTL/PCI-TSM/PCI-IDLE/NS_TNAR )
  );
  X_AND2   \PCI-CNTL/PCI-TSM/PCI-IDLE/$1I496  (
    .I0(\PCI-CNTL/PCI-TSM/PCI-IDLE/EQN-A ),
    .I1(S_DATA_INT),
    .O(\PCI-CNTL/PCI-TSM/PCI-IDLE/DATA_NS_TNAR )
  );
  X_OR2   \PCI-CNTL/PCI-TSM/PCI-IDLE/$1I494  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-IDLE/$1I494/I0 ),
    .I1(\NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-IDLE/$1I494/I1 ),
    .O(\PCI-CNTL/PCI-TSM/PCI-IDLE/$1N483 )
  );
  X_AND2   \PCI-CNTL/PCI-TSM/PCI-IDLE/$1I493  (
    .I0(\PCI-CNTL/PCI-TSM/PCI-IDLE/$1N483 ),
    .I1(\FRAME- ),
    .O(\PCI-CNTL/PCI-TSM/PCI-IDLE/EQN-A )
  );
  X_AND2   \PCI-CNTL/PCI-TSM/PCI-IDLE/$1I369  (
    .I0(\FRAME- ),
    .I1(\PCI-CNTL/PCI-TSM/PCI-IDLE/$1N367 ),
    .O(\PCI-CNTL/PCI-TSM/PCI-IDLE/IDLE_NS_IDLE )
  );
  X_OR2   \PCI-CNTL/PCI-TSM/PCI-IDLE/$1I365  (
    .I0(TURN_AR_INT),
    .I1(IDLE_INT),
    .O(\PCI-CNTL/PCI-TSM/PCI-IDLE/$1N367 )
  );
  X_OR3   \PCI-CNTL/PCI-TSM/PCI-IDLE/$1I337  (
    .I0(\PCI-CNTL/PCI-TSM/PCI-IDLE/BUSY_NS_IDLE ),
    .I1(\PCI-CNTL/PCI-TSM/PCI-IDLE/IDLE_NS_IDLE ),
    .I2(\PCI-CNTL/PCI-TSM/PCI-IDLE/NS_TNAR ),
    .O(\PCI-CNTL/PCI-TSM/PCI-IDLE/NS_IDLE )
  );
  X_AND3   \PCI-CNTL/PCI-TSM/PCI-IDLE/$1I321  (
    .I0(\IRDY- ),
    .I1(\FRAME- ),
    .I2(B_BUSY_INT),
    .O(\PCI-CNTL/PCI-TSM/PCI-IDLE/BUSY_NS_IDLE )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-CNTL/PCI-TSM/PCI-IDLE/IDLE0_FF  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(CLK),
    .I(\PCI-CNTL/PCI-TSM/PCI-IDLE/NS_IDLE ),
    .O(IDLE_INT),
    .RST(GND)
  );
  X_OR4   \PCI-CNTL/PCI-TSM/PCI-BUSY/$1I572  (
    .I0(NlwRenamedSig_OI_BASE_HIT2),
    .I1(NlwRenamedSig_OI_BASE_HIT1),
    .I2(NlwRenamedSig_OI_BASE_HIT0),
    .I3(NlwRenamedSig_OI_CFG_HIT),
    .O(\PCI-CNTL/PCI-TSM/PCI-BUSY/HITIDLEORBUSY )
  );
  X_OR2   \PCI-CNTL/PCI-TSM/PCI-BUSY/$1I547  (
    .I0(\PCI-CNTL/PCI-TSM/PCI-BUSY/BUSY_NS_BUSY ),
    .I1(\PCI-CNTL/PCI-TSM/PCI-BUSY/IDLE_NS_BUSY ),
    .O(\PCI-CNTL/PCI-TSM/PCI-BUSY/NS_BUSY )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-TSM/PCI-BUSY/BUSY_FF  (
    .CE(VCC),
    .CLK(CLK),
    .I(\PCI-CNTL/PCI-TSM/PCI-BUSY/NS_BUSY ),
    .O(B_BUSY_INT),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND2   \PCI-CNTL/PCI-TSM/PCI-BUSY/$1I542  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-BUSY/$1I542/I0 ),
    .I1(\PCI-CNTL/PCI-TSM/PCI-BUSY/EQN-B ),
    .O(\PCI-CNTL/PCI-TSM/PCI-BUSY/BUSY_NS_BUSY )
  );
  X_AND2   \PCI-CNTL/PCI-TSM/PCI-BUSY/$1I521  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-BUSY/$1I521/I0 ),
    .I1(\PCI-CNTL/PCI-TSM/PCI-BUSY/EQN-A ),
    .O(\PCI-CNTL/PCI-TSM/PCI-BUSY/IDLE_NS_BUSY )
  );
  X_OR2   \PCI-CNTL/PCI-TSM/PCI-BUSY/$1I473  (
    .I0(TURN_AR_INT),
    .I1(IDLE_INT),
    .O(\PCI-CNTL/PCI-TSM/PCI-BUSY/$1N476 )
  );
  X_AND2   \PCI-CNTL/PCI-TSM/PCI-BUSY/$1I472  (
    .I0(\PCI-CNTL/PCI-TSM/PCI-BUSY/$1N484 ),
    .I1(B_BUSY_INT),
    .O(\PCI-CNTL/PCI-TSM/PCI-BUSY/EQN-B )
  );
  X_OR2   \PCI-CNTL/PCI-TSM/PCI-BUSY/$1I471  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-BUSY/$1I471/I0 ),
    .I1(\NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-BUSY/$1I471/I1 ),
    .O(\PCI-CNTL/PCI-TSM/PCI-BUSY/$1N484 )
  );
  X_AND2   \PCI-CNTL/PCI-TSM/PCI-BUSY/$1I469  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-BUSY/$1I469/I0 ),
    .I1(\PCI-CNTL/PCI-TSM/PCI-BUSY/$1N476 ),
    .O(\PCI-CNTL/PCI-TSM/PCI-BUSY/EQN-A )
  );
  X_BUF   \PCI-CNTL/PCI-TSM/PCI-BUSY/$1I587/NC  (
    .I(BACKOFF_INT),
    .O(\NLW_PCI-CNTL/PCI-TSM/PCI-BUSY/$1I587/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-CNTL/PCI-TSM/PCI-BUSY/$1I588/NC  (
    .I(S_DATA_INT),
    .O(\NLW_PCI-CNTL/PCI-TSM/PCI-BUSY/$1I588/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-CNTL/PCI-TSM/PCI-BUSY/$1I589/NC  (
    .I(\PCI-CNTL/TSTOP- ),
    .O(\NLW_PCI-CNTL/PCI-TSM/PCI-BUSY/$1I589/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-CNTL/PCI-TSM/PCI-BUSY/$1I590/NC  (
    .I(\PCI-CNTL/TTRDY- ),
    .O(\NLW_PCI-CNTL/PCI-TSM/PCI-BUSY/$1I590/NC_O_UNCONNECTED )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-TSM/PCI-DATA/DATA1_FF  (
    .CE(VCC),
    .CLK(CLK),
    .I(\PCI-CNTL/PCI-TSM/PCI-DATA/NS_DATA ),
    .O(S_DATA),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_OR2   \PCI-CNTL/PCI-TSM/PCI-DATA/$1I670  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-DATA/$1I670/I0 ),
    .I1(\NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-DATA/$1I670/I1 ),
    .O(\PCI-CNTL/PCI-TSM/PCI-DATA/$1N673 )
  );
  X_AND2   \PCI-CNTL/PCI-TSM/PCI-DATA/$1I668  (
    .I0(\PCI-CNTL/PCI-TSM/PCI-DATA/$1N673 ),
    .I1(B_BUSY_INT),
    .O(\PCI-CNTL/PCI-TSM/PCI-DATA/EQN-A )
  );
  X_AND3   \PCI-CNTL/PCI-TSM/PCI-DATA/$1I631  (
    .I0(\PCI-CNTL/PCI-TSM/PCI-DATA/EQN-B ),
    .I1(NlwRenamedSig_OI_CFG_HIT),
    .I2(\PCI-CNTL/PCI-TSM/PCI-DATA/EQN-A ),
    .O(\PCI-CNTL/PCI-TSM/PCI-DATA/CBUSY_NS_DATA )
  );
  X_AND2   \PCI-CNTL/PCI-TSM/PCI-DATA/$1I629  (
    .I0(C_READY),
    .I1(C_TERM),
    .O(\PCI-CNTL/PCI-TSM/PCI-DATA/$1N628 )
  );
  X_OR2   \PCI-CNTL/PCI-TSM/PCI-DATA/$1I627  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-DATA/$1I627/I0 ),
    .I1(\PCI-CNTL/PCI-TSM/PCI-DATA/$1N628 ),
    .O(\PCI-CNTL/PCI-TSM/PCI-DATA/EQN-B )
  );
  X_OR3   \PCI-CNTL/PCI-TSM/PCI-DATA/$1I562  (
    .I0(\PCI-CNTL/PCI-TSM/PCI-DATA/DATA_NS_DATA ),
    .I1(\PCI-CNTL/PCI-TSM/PCI-DATA/BUSY_NS_DATA ),
    .I2(\PCI-CNTL/PCI-TSM/PCI-DATA/CBUSY_NS_DATA ),
    .O(\PCI-CNTL/PCI-TSM/PCI-DATA/NS_DATA )
  );
  X_OR3   \PCI-CNTL/PCI-TSM/PCI-DATA/$1I548  (
    .I0(NlwRenamedSig_OI_BASE_HIT2),
    .I1(NlwRenamedSig_OI_BASE_HIT1),
    .I2(NlwRenamedSig_OI_BASE_HIT0),
    .O(\PCI-CNTL/PCI-TSM/PCI-DATA/HIT )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-TSM/PCI-DATA/DATA0_FF  (
    .CE(VCC),
    .CLK(CLK),
    .I(\PCI-CNTL/PCI-TSM/PCI-DATA/NS_DATA ),
    .O(S_DATA_INT),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND2   \PCI-CNTL/PCI-TSM/PCI-DATA/$1I503  (
    .I0(\PCI-CNTL/PCI-TSM/PCI-DATA/EQN-E ),
    .I1(S_DATA_INT),
    .O(\PCI-CNTL/PCI-TSM/PCI-DATA/DATA_NS_DATA )
  );
  X_AND3   \PCI-CNTL/PCI-TSM/PCI-DATA/$1I482  (
    .I0(\PCI-CNTL/TTRDY- ),
    .I1(\PCI-CNTL/TSTOP- ),
    .I2(\FRAME- ),
    .O(\PCI-CNTL/PCI-TSM/PCI-DATA/$1N495 )
  );
  X_AND2   \PCI-CNTL/PCI-TSM/PCI-DATA/$1I481  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-DATA/$1I481/I0 ),
    .I1(\PCI-CNTL/TSTOP- ),
    .O(\PCI-CNTL/PCI-TSM/PCI-DATA/$1N483 )
  );
  X_AND4   \PCI-CNTL/PCI-TSM/PCI-DATA/$1I480  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-DATA/$1I480/I0 ),
    .I1(\NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-DATA/$1I480/I1 ),
    .I2(\NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-DATA/$1I480/I2 ),
    .I3(\IRDY- ),
    .O(\PCI-CNTL/PCI-TSM/PCI-DATA/$1N497 )
  );
  X_OR3   \PCI-CNTL/PCI-TSM/PCI-DATA/$1I479  (
    .I0(\PCI-CNTL/PCI-TSM/PCI-DATA/$1N495 ),
    .I1(\PCI-CNTL/PCI-TSM/PCI-DATA/$1N483 ),
    .I2(\PCI-CNTL/PCI-TSM/PCI-DATA/$1N497 ),
    .O(\PCI-CNTL/PCI-TSM/PCI-DATA/EQN-E )
  );
  X_AND3   \PCI-CNTL/PCI-TSM/PCI-DATA/$1I465  (
    .I0(\PCI-CNTL/PCI-TSM/PCI-DATA/EQN-D ),
    .I1(\PCI-CNTL/PCI-TSM/PCI-DATA/HIT ),
    .I2(\PCI-CNTL/PCI-TSM/PCI-DATA/EQN-A ),
    .O(\PCI-CNTL/PCI-TSM/PCI-DATA/BUSY_NS_DATA )
  );
  X_OR2   \PCI-CNTL/PCI-TSM/PCI-DATA/$1I453  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-DATA/$1I453/I0 ),
    .I1(\PCI-CNTL/PCI-TSM/PCI-DATA/$1N452 ),
    .O(\PCI-CNTL/PCI-TSM/PCI-DATA/EQN-D )
  );
  X_AND2   \PCI-CNTL/PCI-TSM/PCI-DATA/$1I450  (
    .I0(S_READY),
    .I1(S_TERM),
    .O(\PCI-CNTL/PCI-TSM/PCI-DATA/$1N452 )
  );
  X_BUF   \PCI-CNTL/PCI-TSM/PCI-DATA/$1I568/NC  (
    .I(BACKOFF_INT),
    .O(\NLW_PCI-CNTL/PCI-TSM/PCI-DATA/$1I568/NC_O_UNCONNECTED )
  );
  X_AND2   \PCI-CNTL/PCI-TSM/PCI-BKOF/$1I599  (
    .I0(\PCI-CNTL/PCI-TSM/PCI-BKOF/BKOF_HIT ),
    .I1(\PCI-CNTL/PCI-TSM/PCI-BKOF/EQN-AB ),
    .O(\PCI-CNTL/PCI-TSM/PCI-BKOF/IDLE_BUSY_NS )
  );
  X_OR2   \PCI-CNTL/PCI-TSM/PCI-BKOF/$1I596  (
    .I0(\PCI-CNTL/PCI-TSM/PCI-BKOF/EQN-B ),
    .I1(\PCI-CNTL/PCI-TSM/PCI-BKOF/EQN-A ),
    .O(\PCI-CNTL/PCI-TSM/PCI-BKOF/EQN-AB )
  );
  X_OR2   \PCI-CNTL/PCI-TSM/PCI-BKOF/$1I583  (
    .I0(\PCI-CNTL/PCI-TSM/PCI-BKOF/C_EQN ),
    .I1(\PCI-CNTL/PCI-TSM/PCI-BKOF/S_EQN ),
    .O(\PCI-CNTL/PCI-TSM/PCI-BKOF/BKOF_HIT )
  );
  X_AND3   \PCI-CNTL/PCI-TSM/PCI-BKOF/$1I579  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-BKOF/$1I579/I0 ),
    .I1(S_TERM),
    .I2(\PCI-CNTL/PCI-TSM/PCI-BKOF/HIT ),
    .O(\PCI-CNTL/PCI-TSM/PCI-BKOF/S_EQN )
  );
  X_AND3   \PCI-CNTL/PCI-TSM/PCI-BKOF/$1I575  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-BKOF/$1I575/I0 ),
    .I1(C_TERM),
    .I2(NlwRenamedSig_OI_CFG_HIT),
    .O(\PCI-CNTL/PCI-TSM/PCI-BKOF/C_EQN )
  );
  X_OR2   \PCI-CNTL/PCI-TSM/PCI-BKOF/$1I526  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-BKOF/$1I526/I0 ),
    .I1(\NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-BKOF/$1I526/I1 ),
    .O(\PCI-CNTL/PCI-TSM/PCI-BKOF/$1N531 )
  );
  X_AND2   \PCI-CNTL/PCI-TSM/PCI-BKOF/$1I525  (
    .I0(\PCI-CNTL/PCI-TSM/PCI-BKOF/$1N531 ),
    .I1(B_BUSY_INT),
    .O(\PCI-CNTL/PCI-TSM/PCI-BKOF/EQN-B )
  );
  X_OR2   \PCI-CNTL/PCI-TSM/PCI-BKOF/$1I508  (
    .I0(\PCI-CNTL/PCI-TSM/PCI-BKOF/DATA_NS ),
    .I1(\PCI-CNTL/PCI-TSM/PCI-BKOF/IDLE_BUSY_NS ),
    .O(\PCI-CNTL/PCI-TSM/PCI-BKOF/NS_BKOF )
  );
  X_OR3   \PCI-CNTL/PCI-TSM/PCI-BKOF/$1I492  (
    .I0(NlwRenamedSig_OI_BASE_HIT2),
    .I1(NlwRenamedSig_OI_BASE_HIT1),
    .I2(NlwRenamedSig_OI_BASE_HIT0),
    .O(\PCI-CNTL/PCI-TSM/PCI-BKOF/HIT )
  );
  X_AND2   \PCI-CNTL/PCI-TSM/PCI-BKOF/$1I486  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-BKOF/$1I486/I0 ),
    .I1(BACKOFF_INT),
    .O(\PCI-CNTL/PCI-TSM/PCI-BKOF/BKOF_NS_BKOF )
  );
  X_AND2   \PCI-CNTL/PCI-TSM/PCI-BKOF/$1I481  (
    .I0(\PCI-CNTL/PCI-TSM/PCI-BKOF/EQN-E ),
    .I1(S_DATA_INT),
    .O(\PCI-CNTL/PCI-TSM/PCI-BKOF/DATA_NS_BKOF )
  );
  X_AND2   \PCI-CNTL/PCI-TSM/PCI-BKOF/$1I476  (
    .I0(\PCI-CNTL/PCI-TSM/PCI-BKOF/$1N479 ),
    .I1(\PCI-CNTL/PCI-TSM/PCI-BKOF/$1N477 ),
    .O(\PCI-CNTL/PCI-TSM/PCI-BKOF/EQN-E )
  );
  X_OR2   \PCI-CNTL/PCI-TSM/PCI-BKOF/$1I475  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-BKOF/$1I475/I0 ),
    .I1(\PCI-CNTL/TTRDY- ),
    .O(\PCI-CNTL/PCI-TSM/PCI-BKOF/$1N479 )
  );
  X_AND2   \PCI-CNTL/PCI-TSM/PCI-BKOF/$1I474  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-BKOF/$1I474/I0 ),
    .I1(\NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-BKOF/$1I474/I1 ),
    .O(\PCI-CNTL/PCI-TSM/PCI-BKOF/$1N477 )
  );
  X_OR2   \PCI-CNTL/PCI-TSM/PCI-BKOF/$1I460  (
    .I0(TURN_AR_INT),
    .I1(IDLE_INT),
    .O(\PCI-CNTL/PCI-TSM/PCI-BKOF/TURNIDLE )
  );
  X_AND2   \PCI-CNTL/PCI-TSM/PCI-BKOF/$1I458  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-BKOF/$1I458/I0 ),
    .I1(\PCI-CNTL/PCI-TSM/PCI-BKOF/TURNIDLE ),
    .O(\PCI-CNTL/PCI-TSM/PCI-BKOF/EQN-A )
  );
  X_OR2   \PCI-CNTL/PCI-TSM/PCI-BKOF/$1I400  (
    .I0(\PCI-CNTL/PCI-TSM/PCI-BKOF/BKOF_NS_BKOF ),
    .I1(\PCI-CNTL/PCI-TSM/PCI-BKOF/DATA_NS_BKOF ),
    .O(\PCI-CNTL/PCI-TSM/PCI-BKOF/DATA_NS )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-TSM/PCI-BKOF/BKOF_FF  (
    .CE(VCC),
    .CLK(CLK),
    .I(\PCI-CNTL/PCI-TSM/PCI-BKOF/NS_BKOF ),
    .O(BACKOFF_INT),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_ZERO   \PCI-CNTL/PCI-TSM/$1I426/$1I2218  (
    .O(\PCI-CNTL/PCI-TSM/$1I426/$1N2216 )
  );
  X_BUF   \PCI-CNTL/PCI-TSM/$1I426/L  (
    .I(\PCI-CNTL/PCI-TSM/$1I426/$1N2216 ),
    .O(TURN_AR_INT)
  );
  X_BUF   \PCI-CNTL/PCI-TSM/$1I489/NC  (
    .I(\PCI-CNTL/S_ABORT ),
    .O(\NLW_PCI-CNTL/PCI-TSM/$1I489/NC_O_UNCONNECTED )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/$1I1430  (
    .I0(\PCI-CNTL/PCI-OFCN/$1N1433 ),
    .I1(\PCI-CNTL/PCI-OFCN/$1N1431 ),
    .O(\PCI-CNTL/PCI-OFCN/NL_MEM )
  );
  X_OR4   \PCI-CNTL/PCI-OFCN/$1I1429  (
    .I0(NL_MEM0),
    .I1(NL_MEM1),
    .I2(NL_MEM2),
    .I3(NL_MEM3),
    .O(\PCI-CNTL/PCI-OFCN/$1N1433 )
  );
  X_OR4   \PCI-CNTL/PCI-OFCN/$1I1428  (
    .I0(NL_MEM4),
    .I1(NL_MEM5),
    .I2(NL_MEM6),
    .I3(NL_MEM7),
    .O(\PCI-CNTL/PCI-OFCN/$1N1431 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-CNTL/PCI-OFCN/PCI-AK64/ACK64  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(ACK64_CE),
    .CLK(CLK),
    .I(\NS_ACK64- ),
    .O(\TACK64_I- ),
    .RST(GND)
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-AK64/$3I855  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-AK64/NS_HIT ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-AK64/$3N836 ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-AK64/$3I855/O )
  );
  X_MUX2   \PCI-CNTL/PCI-OFCN/PCI-AK64/$3I848  (
    .IA(\PCI-CNTL/PCI-OFCN/PCI-AK64/NS_F0 ),
    .IB(\PCI-CNTL/PCI-OFCN/PCI-AK64/NS_F1 ),
    .O(\NS_ACK64- ),
    .SEL(REQ64_I)
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-CNTL/PCI-OFCN/PCI-AK64/ACK64Q-  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(CLK),
    .I(\TACK64_I- ),
    .O(\PCI-CNTL/TACK64- ),
    .RST(GND)
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-AK64/$2I977  (
    .I0(\PCI-CNTL/TSTOP- ),
    .I1(\PCI-CNTL/TTRDY- ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-AK64/$2N962 )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-AK64/$2I975  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-AK64/BKOF_NS_BKOF ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-AK64/DATA_NS_DATA_OR_BKOF1 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-AK64/$2N974 )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-AK64/$2I973  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-AK64/$2N970 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-AK64/EQN-C ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-AK64/NS_F0_I1 )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-AK64/$2I972  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-AK64/$2N969 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-AK64/EQN-C ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-AK64/NS_F0_I0 )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-AK64/$2I971  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-AK64/$2I971/I0 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-AK64/$2N968 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-AK64/$2N969 )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-AK64/$2I965  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-AK64/$2I965/I0 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-AK64/$2N974 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-AK64/$2N970 )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-AK64/$2I964  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-AK64/BKOF_NS_BKOF ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-AK64/DATA_NS_DATA_OR_BKOF0 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-AK64/$2N968 )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-AK64/$2I959  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-AK64/$2N982 ),
    .I1(S_DATA_INT),
    .O(\PCI-CNTL/PCI-OFCN/PCI-AK64/DATA_NS_DATA_OR_BKOF0 )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-AK64/$2I958  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-AK64/$2I958/I0 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-AK64/$2N962 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-AK64/$2N982 )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-AK64/$2I951  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-AK64/$2I951/I0 ),
    .I1(BACKOFF_INT),
    .O(\PCI-CNTL/PCI-OFCN/PCI-AK64/BKOF_NS_BKOF )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-AK64/$2I948  (
    .I0(\TTRDY_I- ),
    .I1(\PCI-CNTL/S_ABORT ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-AK64/DUCKLING )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-AK64/$2I941  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-AK64/$2I941/I0 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-AK64/$2N937 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-AK64/$2N931 )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-AK64/$2I940  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-AK64/$2N931 ),
    .I1(S_DATA_INT),
    .O(\PCI-CNTL/PCI-OFCN/PCI-AK64/DATA_NS_DATA_OR_BKOF1 )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-AK64/$2I936  (
    .I0(\PCI-CNTL/TSTOP- ),
    .I1(\PCI-CNTL/TTRDY- ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-AK64/$2N937 )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-AK64/$1I837  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-AK64/$1I837/I0 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-AK64/$1N809 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-AK64/EQN-F1A )
  );
  X_OR3   \PCI-CNTL/PCI-OFCN/PCI-AK64/$1I831  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-AK64/EQN-F1A ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-AK64/EQN-C ),
    .I2(\PCI-CNTL/PCI-OFCN/PCI-AK64/NS_HIT ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-AK64/$1N801 )
  );
  X_AND3   \PCI-CNTL/PCI-OFCN/PCI-AK64/$1I830  (
    .I0(\TTRDY_I- ),
    .I1(\PCI-CNTL/TSTOP- ),
    .I2(\TSTOP_I- ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-AK64/LATE_GATE )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-AK64/$1I808  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-AK64/$1N846 ),
    .I1(\PCI-CNTL/PCI-OFCN/ACKHIT ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-AK64/EQN-C )
  );
  X_OR3   \PCI-CNTL/PCI-OFCN/PCI-AK64/$1I807  (
    .I0(BH64_2),
    .I1(BH64_1),
    .I2(BH64_0),
    .O(\PCI-CNTL/PCI-OFCN/ACKHIT )
  );
  X_OR3   \PCI-CNTL/PCI-OFCN/PCI-AK64/$1I806  (
    .I0(NS_BH64_2),
    .I1(NS_BH64_1),
    .I2(NS_BH64_0),
    .O(\PCI-CNTL/PCI-OFCN/PCI-AK64/NS_HIT )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-AK64/$1I797  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-AK64/$1I797/I0 ),
    .I1(BACKOFF_INT),
    .O(\PCI-CNTL/PCI-OFCN/PCI-AK64/$1N794 )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-AK64/$1I796  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-AK64/$1I796/I0 ),
    .I1(\PCI-CNTL/TTRDY- ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-AK64/$1N789 )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-AK64/$1I791  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-AK64/$1N794 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-AK64/$1N795 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-AK64/$1N809 )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-AK64/$1I790  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-AK64/$1N789 ),
    .I1(S_DATA_INT),
    .O(\PCI-CNTL/PCI-OFCN/PCI-AK64/$1N795 )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-AK64/$1I787  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-AK64/$1N801 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-AK64/LATE_GATE ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-AK64/$1I787/O )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-AK64/$1I781  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-AK64/$1I781/I0 ),
    .I1(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-AK64/$1I781/I1 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-AK64/$1N782 )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-AK64/$1I780  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-AK64/$1N782 ),
    .I1(B_BUSY_INT),
    .O(\PCI-CNTL/PCI-OFCN/PCI-AK64/$1N846 )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-AK64/$3I854/$1I9  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-AK64/NS_F0_I1 ),
    .I1(IRDY_M),
    .O(\PCI-CNTL/PCI-OFCN/PCI-AK64/$3I854/M1 )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-AK64/$3I854/$1I8  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-AK64/$3I854/M1 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-AK64/$3I854/M0 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-AK64/$3N836 )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-AK64/$3I854/$1I7  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-AK64/$3I854/$1I7/I0 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-AK64/NS_F0_I0 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-AK64/$3I854/M0 )
  );
  X_ONE   \PCI-CNTL/PCI-OFCN/PCI-AK64/$3I864/$1I2220  (
    .O(\PCI-CNTL/PCI-OFCN/PCI-AK64/$3I864/$1N2216 )
  );
  X_BUF   \PCI-CNTL/PCI-OFCN/PCI-AK64/$3I864/H  (
    .I(\PCI-CNTL/PCI-OFCN/PCI-AK64/$3I864/$1N2216 ),
    .O(ACK64_CE)
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-DSEL/$3I795  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-DSEL/NS_HIT ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-DSEL/$3N806 ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-DSEL/$3I795/O )
  );
  X_MUX2   \PCI-CNTL/PCI-OFCN/PCI-DSEL/$3I781  (
    .IA(\PCI-CNTL/PCI-OFCN/PCI-DSEL/NS_F0 ),
    .IB(\PCI-CNTL/PCI-OFCN/PCI-DSEL/NS_F1 ),
    .O(\NS_DEVSEL- ),
    .SEL(FRAME_I)
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-CNTL/PCI-OFCN/PCI-DSEL/DEVSEL  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(DEVSEL_CE),
    .CLK(CLK),
    .I(\NS_DEVSEL- ),
    .O(\TDEVSEL_I- ),
    .RST(GND)
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-CNTL/PCI-OFCN/PCI-DSEL/DEVSELQ-  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(CLK),
    .I(\TDEVSEL_I- ),
    .O(\PCI-CNTL/TDEVSEL- ),
    .RST(GND)
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-DSEL/$2I983  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-DSEL/$2I983/I0 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-DSEL/$2N979 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-DSEL/$2N972 )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-DSEL/$2I982  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-DSEL/$2N972 ),
    .I1(S_DATA_INT),
    .O(\PCI-CNTL/PCI-OFCN/PCI-DSEL/DATA_NS_DATA_OR_BKOF1 )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-DSEL/$2I977  (
    .I0(\PCI-CNTL/TSTOP- ),
    .I1(\PCI-CNTL/TTRDY- ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-DSEL/$2N979 )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-DSEL/$2I959  (
    .I0(\TTRDY_I- ),
    .I1(\PCI-CNTL/S_ABORT ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-DSEL/DUCKLING )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-DSEL/$2I951  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-DSEL/$2I951/I0 ),
    .I1(BACKOFF_INT),
    .O(\PCI-CNTL/PCI-OFCN/PCI-DSEL/BKOF_NS_BKOF )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-DSEL/$2I933  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-DSEL/$2N938 ),
    .I1(S_DATA_INT),
    .O(\PCI-CNTL/PCI-OFCN/PCI-DSEL/DATA_NS_DATA_OR_BKOF0 )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-DSEL/$2I932  (
    .I0(\PCI-CNTL/TSTOP- ),
    .I1(\PCI-CNTL/TTRDY- ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-DSEL/$2N939 )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-DSEL/$2I931  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-DSEL/$2I931/I0 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-DSEL/$2N939 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-DSEL/$2N938 )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-DSEL/$2I914  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-DSEL/$2I914/I0 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-DSEL/$2N899 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-DSEL/$2N917 )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-DSEL/$2I909  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-DSEL/BKOF_NS_BKOF ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-DSEL/DATA_NS_DATA_OR_BKOF0 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-DSEL/$2N899 )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-DSEL/$2I897  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-DSEL/$2N917 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-DSEL/EQN-C ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-DSEL/NS_F0_I0 )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-DSEL/$2I896  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-DSEL/$2N875 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-DSEL/EQN-C ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-DSEL/NS_F0_I1 )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-DSEL/$2I883  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-DSEL/BKOF_NS_BKOF ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-DSEL/DATA_NS_DATA_OR_BKOF1 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-DSEL/$2N893 )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-DSEL/$2I878  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-DSEL/$2I878/I0 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-DSEL/$2N893 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-DSEL/$2N875 )
  );
  X_AND3   \PCI-CNTL/PCI-OFCN/PCI-DSEL/$1I927  (
    .I0(\TTRDY_I- ),
    .I1(\PCI-CNTL/TSTOP- ),
    .I2(\TSTOP_I- ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-DSEL/LATE_GATE )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-DSEL/$1I801  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-DSEL/$1N919 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-DSEL/LATE_GATE ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-DSEL/$1I801/O )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-DSEL/$1I769  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-DSEL/$1N783 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-DSEL/$1N784 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-DSEL/$1N790 )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-DSEL/$1I768  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-DSEL/$1I768/I0 ),
    .I1(\PCI-CNTL/TTRDY- ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-DSEL/$1N923 )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-DSEL/$1I766  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-DSEL/$1N923 ),
    .I1(S_DATA_INT),
    .O(\PCI-CNTL/PCI-OFCN/PCI-DSEL/$1N784 )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-DSEL/$1I760  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-DSEL/$1I760/I0 ),
    .I1(BACKOFF_INT),
    .O(\PCI-CNTL/PCI-OFCN/PCI-DSEL/$1N783 )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-DSEL/$1I758  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-DSEL/$1I758/I0 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-DSEL/$1N790 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-DSEL/EQN-F1A )
  );
  X_OR3   \PCI-CNTL/PCI-OFCN/PCI-DSEL/$1I1035  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-DSEL/EQN-F1A ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-DSEL/EQN-C ),
    .I2(\PCI-CNTL/PCI-OFCN/PCI-DSEL/NS_HIT ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-DSEL/$1N919 )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-DSEL/$1I1034  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-DSEL/$1N1033 ),
    .I1(\PCI-CNTL/PCI-OFCN/HIT ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-DSEL/EQN-C )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-DSEL/$1I1028  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-DSEL/$1I1028/I0 ),
    .I1(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-DSEL/$1I1028/I1 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-DSEL/$1N1030 )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-DSEL/$1I1027  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-DSEL/$1N1030 ),
    .I1(B_BUSY_INT),
    .O(\PCI-CNTL/PCI-OFCN/PCI-DSEL/$1N1033 )
  );
  X_OR4   \PCI-CNTL/PCI-OFCN/PCI-DSEL/$1I1022  (
    .I0(NlwRenamedSig_OI_CFG_HIT),
    .I1(NlwRenamedSig_OI_BASE_HIT2),
    .I2(NlwRenamedSig_OI_BASE_HIT1),
    .I3(NlwRenamedSig_OI_BASE_HIT0),
    .O(\PCI-CNTL/PCI-OFCN/HIT )
  );
  X_OR4   \PCI-CNTL/PCI-OFCN/PCI-DSEL/$1I1015  (
    .I0(\PCI-CNTL/NS_CFG_HIT ),
    .I1(NS_BASE_HIT2),
    .I2(NS_BASE_HIT1),
    .I3(NS_BASE_HIT0),
    .O(\PCI-CNTL/PCI-OFCN/PCI-DSEL/NS_HIT )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-DSEL/$3I798/$1I9  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-DSEL/NS_F0_I1 ),
    .I1(IRDY_M),
    .O(\PCI-CNTL/PCI-OFCN/PCI-DSEL/$3I798/M1 )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-DSEL/$3I798/$1I8  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-DSEL/$3I798/M1 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-DSEL/$3I798/M0 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-DSEL/$3N806 )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-DSEL/$3I798/$1I7  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-DSEL/$3I798/$1I7/I0 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-DSEL/NS_F0_I0 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-DSEL/$3I798/M0 )
  );
  X_ONE   \PCI-CNTL/PCI-OFCN/PCI-DSEL/$3I813/$1I2220  (
    .O(\PCI-CNTL/PCI-OFCN/PCI-DSEL/$3I813/$1N2216 )
  );
  X_BUF   \PCI-CNTL/PCI-OFCN/PCI-DSEL/$3I813/H  (
    .I(\PCI-CNTL/PCI-OFCN/PCI-DSEL/$3I813/$1N2216 ),
    .O(DEVSEL_CE)
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-CNTL/PCI-OFCN/PCI-TRDY/S1FF  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(CLK),
    .I(\PCI-CNTL/PCI-OFCN/PCI-TRDY/S_FIRSTIN ),
    .O(S_FIRST),
    .RST(GND)
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-TRDY/$4I977  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$4I977/I0 ),
    .I1(\TTRDY_I- ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-TRDY/$4N968 )
  );
  X_MUX2   \PCI-CNTL/PCI-OFCN/PCI-TRDY/$4I962  (
    .IA(\PCI-CNTL/PCI-OFCN/PCI-TRDY/S_FIRST0 ),
    .IB(\PCI-CNTL/PCI-OFCN/PCI-TRDY/S_FIRST1 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-TRDY/S_FIRSTIN ),
    .SEL(FRAME_I)
  );
  X_AND3   \PCI-CNTL/PCI-OFCN/PCI-TRDY/$4I1063  (
    .I0(S_FIRST),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-TRDY/SWAN0 ),
    .I2(\PCI-CNTL/PCI-OFCN/PCI-TRDY/$4N968 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-TRDY/SF0_I1 )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-TRDY/$4I1057  (
    .I0(S_FIRST),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-TRDY/$4N1042 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-TRDY/SF0_I0 )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-TRDY/$4I1044  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$4I1044/I0 ),
    .I1(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$4I1044/I1 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-TRDY/$4N1052 )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-TRDY/$4I1043  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-TRDY/$4N1052 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-TRDY/SWAN0 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-TRDY/$4N1042 )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-TRDY/$4I1029  (
    .I0(IDLE_INT),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-TRDY/$4N1030 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-TRDY/S_FIRST0 )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-TRDY/$4I1010  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$4I1010/I0 ),
    .I1(\TTRDY_I- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$4I1010/O )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-TRDY/$4I1005  (
    .I0(S_FIRST),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-TRDY/$4N1002 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-TRDY/$4N1008 )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-TRDY/$4I1004  (
    .I0(IDLE_INT),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-TRDY/$4N1008 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-TRDY/S_FIRST1 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-CNTL/PCI-OFCN/PCI-TRDY/TRDY  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(TRDY_CE),
    .CLK(CLK),
    .I(\NS_TRDY- ),
    .O(\TTRDY_I- ),
    .RST(GND)
  );
  X_MUX2   \PCI-CNTL/PCI-OFCN/PCI-TRDY/$3I928  (
    .IA(\PCI-CNTL/PCI-OFCN/PCI-TRDY/SWAN1 ),
    .IB(\PCI-CNTL/PCI-OFCN/PCI-TRDY/SWAN2 ),
    .O(\NS_TRDY- ),
    .SEL(FRAME_I)
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-CNTL/PCI-OFCN/PCI-TRDY/TRDYQ  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(CLK),
    .I(\TTRDY_I- ),
    .O(\PCI-CNTL/TTRDY- ),
    .RST(GND)
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-TRDY/$3I856  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$3I856/I0 ),
    .I1(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$3I856/I1 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-TRDY/TRDY_OFF )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-TRDY/$3I825  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$3I825/I0 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-TRDY/TRDY_OFF ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-TRDY/$3N837 )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-TRDY/$3I823  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$3I823/I0 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-TRDY/SWAN0 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-TRDY/$3N833 )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-TRDY/$3I822  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$3I822/I0 ),
    .I1(\TTRDY_I- ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-TRDY/HOLD_TRDY )
  );
  X_OR3   \PCI-CNTL/PCI-OFCN/PCI-TRDY/$3I821  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-TRDY/$3N837 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-TRDY/$3N833 ),
    .I2(\PCI-CNTL/PCI-OFCN/PCI-TRDY/$3N835 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-TRDY/SWAN1 )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-TRDY/$3I820  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-TRDY/SWAN0 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-TRDY/HOLD_TRDY ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-TRDY/$3N835 )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-TRDY/$3I616  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$3I616/I0 ),
    .I1(\TTRDY_I- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$3I616/O )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I785  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I785/I0 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-TRDY/$1N786 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-TRDY/EQN-F )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I768  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I768/I0 ),
    .I1(\TDEVSEL_I- ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-TRDY/$1N763 )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I767  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-TRDY/NS_TRDY- ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-TRDY/$1N763 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-TRDY/SWAN0 )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I746  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-TRDY/DATA_NS_DATA ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-TRDY/CRABILL ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I746/O )
  );
  X_AND3   \PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I745  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-TRDY/EQN-F ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-TRDY/BUSY_NS_DATA ),
    .I2(\PCI-CNTL/PCI-OFCN/PCI-TRDY/EQN-A ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-TRDY/CRABILL )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I742  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-TRDY/C_EQN ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-TRDY/S_EQN ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-TRDY/BUSY_NS_DATA )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I736  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-TRDY/$1N738 ),
    .I1(NlwRenamedSig_OI_CFG_HIT),
    .O(\PCI-CNTL/PCI-OFCN/PCI-TRDY/C_EQN )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I732  (
    .I0(C_READY),
    .I1(C_TERM),
    .O(\PCI-CNTL/PCI-OFCN/PCI-TRDY/$1N735 )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I731  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I731/I0 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-TRDY/$1N735 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-TRDY/$1N738 )
  );
  X_OR3   \PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I724  (
    .I0(NlwRenamedSig_OI_BASE_HIT2),
    .I1(NlwRenamedSig_OI_BASE_HIT1),
    .I2(NlwRenamedSig_OI_BASE_HIT0),
    .O(\PCI-CNTL/PCI-OFCN/PCI-TRDY/HIT )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I723  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-TRDY/EQN-D ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-TRDY/HIT ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-TRDY/S_EQN )
  );
  X_AND3   \PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I705  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-TRDY/$1N466 ),
    .I1(NlwRenamedSig_OI_S_WRDN),
    .I2(B_BUSY_INT),
    .O(\PCI-CNTL/PCI-OFCN/PCI-TRDY/EQN-A )
  );
  X_AND3   \PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I503  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-TRDY/EQN-F ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-TRDY/EQN-E ),
    .I2(S_DATA_INT),
    .O(\PCI-CNTL/PCI-OFCN/PCI-TRDY/DATA_NS_DATA )
  );
  X_AND3   \PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I482  (
    .I0(\PCI-CNTL/TTRDY- ),
    .I1(\PCI-CNTL/TSTOP- ),
    .I2(\FRAME- ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-TRDY/$1N495 )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I481  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I481/I0 ),
    .I1(\PCI-CNTL/TSTOP- ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-TRDY/$1N637 )
  );
  X_AND4   \PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I480  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I480/I0 ),
    .I1(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I480/I1 ),
    .I2(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I480/I2 ),
    .I3(\IRDY- ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-TRDY/$1N497 )
  );
  X_OR3   \PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I479  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-TRDY/$1N495 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-TRDY/$1N637 ),
    .I2(\PCI-CNTL/PCI-OFCN/PCI-TRDY/$1N497 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-TRDY/EQN-E )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I459  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I459/I0 ),
    .I1(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I459/I1 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-TRDY/$1N466 )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I453  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I453/I0 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-TRDY/$1N452 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-TRDY/EQN-D )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I450  (
    .I0(S_READY),
    .I1(S_TERM),
    .O(\PCI-CNTL/PCI-OFCN/PCI-TRDY/$1N452 )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I782/$1I9  (
    .I0(C_READY),
    .I1(\PCI-CNTL/CFG_CYC ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I782/M1 )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I782/$1I8  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I782/M1 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I782/M0 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-TRDY/$1N786 )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I782/$1I7  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I782/$1I7/I0 ),
    .I1(S_READY),
    .O(\PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I782/M0 )
  );
  X_ONE   \PCI-CNTL/PCI-OFCN/PCI-TRDY/$3I957/$1I2220  (
    .O(\PCI-CNTL/PCI-OFCN/PCI-TRDY/$3I957/$1N2216 )
  );
  X_BUF   \PCI-CNTL/PCI-OFCN/PCI-TRDY/$3I957/H  (
    .I(\PCI-CNTL/PCI-OFCN/PCI-TRDY/$3I957/$1N2216 ),
    .O(TRDY_CE)
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-TRDY/$4I1028/$1I9  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-TRDY/SF0_I1 ),
    .I1(IRDY_M),
    .O(\PCI-CNTL/PCI-OFCN/PCI-TRDY/$4I1028/M1 )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-TRDY/$4I1028/$1I8  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-TRDY/$4I1028/M1 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-TRDY/$4I1028/M0 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-TRDY/$4N1030 )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-TRDY/$4I1028/$1I7  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$4I1028/$1I7/I0 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-TRDY/SF0_I0 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-TRDY/$4I1028/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-CNTL/PCI-OFCN/PCI-STOP/STOPQ  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(CLK),
    .I(\TSTOP_I- ),
    .O(\PCI-CNTL/TSTOP- ),
    .RST(GND)
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-CNTL/PCI-OFCN/PCI-STOP/STOP  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(STOP_CE),
    .CLK(CLK),
    .I(\NS_STOP- ),
    .O(\TSTOP_I- ),
    .RST(GND)
  );
  X_MUX2   \PCI-CNTL/PCI-OFCN/PCI-STOP/$3I1328  (
    .IA(\PCI-CNTL/PCI-OFCN/PCI-STOP/NS_0 ),
    .IB(\PCI-CNTL/PCI-OFCN/PCI-STOP/NS_1 ),
    .O(\NS_STOP- ),
    .SEL(IRDY_M)
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-STOP/$3I1287  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$3I1287/I0 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-STOP/$3N1288 ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$3I1287/O )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-STOP/$3I1286  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$3I1286/I0 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-STOP/$3N1277 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-STOP/$3N1288 )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-STOP/$3I1284  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$3I1284/I0 ),
    .I1(FRAME_I),
    .O(\PCI-CNTL/PCI-OFCN/PCI-STOP/$3N1280 )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-STOP/$3I1276  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-STOP/SUB_DATA ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-STOP/PRE_DATA ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-STOP/$3N1277 )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-STOP/$3I1263  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$3I1263/I0 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-STOP/PRE_NS ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$3I1263/O )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-STOP/$3I1261  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-STOP/$3N1257 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-STOP/$3N1259 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-STOP/$3N1256 )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-STOP/$3I1260  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$3I1260/I0 ),
    .I1(FRAME_I),
    .O(\PCI-CNTL/PCI-OFCN/PCI-STOP/$3N1259 )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-STOP/$3I1258  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$3I1258/I0 ),
    .I1(FRAME_I),
    .O(\PCI-CNTL/PCI-OFCN/PCI-STOP/$3N1257 )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1504  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1504/I0 ),
    .I1(\PCI-CNTL/TSTOP- ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-STOP/NUPUR )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1502  (
    .I0(\PCI-CNTL/TDEVSEL- ),
    .I1(\TDEVSEL_I- ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-STOP/$1N1503 )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1495  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-STOP/$1N1500 ),
    .I1(\PCI-CNTL/S_ABORT ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-STOP/JAYANT )
  );
  X_AND3   \PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1480  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1480/I0 ),
    .I1(\TTRDY_I- ),
    .I2(\PCI-CNTL/PCI-OFCN/PCI-STOP/NUPUR ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-STOP/IDATA_WIN )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1456  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-STOP/NUPUR ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-STOP/JAYANT ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-STOP/$1N1459 )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1454  (
    .I0(\TTRDY_I- ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-STOP/$1N1459 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-STOP/SUB_DATA )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1451  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-STOP/$1N1159 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-STOP/PRE_DATA ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-STOP/$1N1453 )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1450  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1450/I0 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-STOP/$1N1453 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-STOP/PRE_NS )
  );
  X_INV   \PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1440  (
    .I(\TTRDY_I- ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-STOP/$1N1434 )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1439  (
    .I0(B_BUSY_INT),
    .I1(IDLE_INT),
    .O(\PCI-CNTL/PCI-OFCN/PCI-STOP/$1N1438 )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1417  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-STOP/TERM ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-STOP/TERM_OTHER ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-STOP/TERMINATE )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1415  (
    .I0(\PCI-CNTL/S_ABORT ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-STOP/DIS_WDATA ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-STOP/TERM_OTHER )
  );
  X_OR4   \PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1360  (
    .I0(NlwRenamedSig_OI_CFG_HIT),
    .I1(NlwRenamedSig_OI_BASE_HIT2),
    .I2(NlwRenamedSig_OI_BASE_HIT1),
    .I3(NlwRenamedSig_OI_BASE_HIT0),
    .O(\PCI-CNTL/PCI-OFCN/PCI-STOP/HIT )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1292  (
    .I0(S_READY),
    .I1(\PCI-CNTL/PCI-OFCN/NL_MEM ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-STOP/DIS_WDATA )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1253  (
    .I0(B_BUSY_INT),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-STOP/HIT ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-STOP/PRE_DEVSEL )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1252  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-STOP/TERMINATE ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-STOP/$1N1266 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-STOP/PRE_DATA )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1251  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-STOP/IDATA_WIN ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-STOP/FAST_TERM_WIN ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-STOP/$1N1266 )
  );
  X_AND3   \PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1248  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1248/I0 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-STOP/WR_OR_NRDY ),
    .I2(\PCI-CNTL/PCI-OFCN/PCI-STOP/PRE_DEVSEL ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-STOP/FAST_TERM_WIN )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1182  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-STOP/NUPUR ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-STOP/JAYANT ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-STOP/$1N1159 )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1060  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1060/I0 ),
    .I1(NlwRenamedSig_OI_S_WRDN),
    .O(\PCI-CNTL/PCI-OFCN/PCI-STOP/WR_OR_NRDY )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1368/$1I9  (
    .I0(C_TERM),
    .I1(\PCI-CNTL/CFG_CYC ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1368/M1 )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1368/$1I8  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1368/M1 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1368/M0 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-STOP/TERM )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1368/$1I7  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1368/$1I7/I0 ),
    .I1(S_TERM),
    .O(\PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1368/M0 )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1373/$1I9  (
    .I0(C_READY),
    .I1(\PCI-CNTL/CFG_CYC ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1373/M1 )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1373/$1I8  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1373/M1 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1373/M0 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-STOP/READY )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1373/$1I7  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1373/$1I7/I0 ),
    .I1(S_READY),
    .O(\PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1373/M0 )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1437/$1I2214  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-STOP/$1N1434 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-STOP/I_DATA_FLAG ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1437/$1N2215 )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1437/$1I2213  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1437/$1I2213/I0 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1437/$1N2215 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1437/D )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1437/FDCE  (
    .CE(VCC),
    .CLK(CLK),
    .I(\PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1437/D ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-STOP/I_DATA_FLAG ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1499/$1I9  (
    .I0(C_TERM),
    .I1(\PCI-CNTL/CFG_CYC ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1499/M1 )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1499/$1I8  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1499/M1 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1499/M0 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-STOP/$1N1500 )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1499/$1I7  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1499/$1I7/I0 ),
    .I1(S_TERM),
    .O(\PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1499/M0 )
  );
  X_ONE   \PCI-CNTL/PCI-OFCN/PCI-STOP/$3I1332/$1I2220  (
    .O(\PCI-CNTL/PCI-OFCN/PCI-STOP/$3I1332/$1N2216 )
  );
  X_BUF   \PCI-CNTL/PCI-OFCN/PCI-STOP/$3I1332/H  (
    .I(\PCI-CNTL/PCI-OFCN/PCI-STOP/$3I1332/$1N2216 ),
    .O(STOP_CE)
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-XOE/$6I996  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-XOE/SET_B64 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-XOE/END64 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/NS-OE_ADO_B64 )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-XOE/$6I971  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-XOE/SET_LB64 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-XOE/END64 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/NS-OE_ADO_LB64 )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-XOE/$6I970  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$6I970/I0 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-XOE/BEGIN64 ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$6I970/O )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-XOE/$6I969  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$6I969/I0 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-XOE/BEGIN64 ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$6I969/O )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-XOE/$6I968  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-XOE/SET_LT64 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-XOE/END64 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/NS-OE_ADO_LT64 )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-XOE/$6I967  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-XOE/SET_T64 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-XOE/END64 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/NS-OE_ADO_T64 )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-XOE/$6I966  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$6I966/I0 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-XOE/BEGIN64 ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$6I966/O )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-XOE/$6I965  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$6I965/I0 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-XOE/BEGIN64 ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$6I965/O )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-CNTL/PCI-OFCN/PCI-XOE/OE_ADO_B64  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(CLK),
    .I(\PCI-CNTL/PCI-OFCN/PCI-XOE/NS-OE_ADO_B64 ),
    .O(OE_AD_T_B64),
    .RST(GND)
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-CNTL/PCI-OFCN/PCI-XOE/OE_ADO_LT64  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(CLK),
    .I(\PCI-CNTL/PCI-OFCN/PCI-XOE/NS-OE_ADO_LT64 ),
    .O(OE_AD_T_LT64),
    .RST(GND)
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-CNTL/PCI-OFCN/PCI-XOE/OE_ADO_LB64  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(CLK),
    .I(\PCI-CNTL/PCI-OFCN/PCI-XOE/NS-OE_ADO_LB64 ),
    .O(OE_AD_T_LB64),
    .RST(GND)
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-CNTL/PCI-OFCN/PCI-XOE/OE_ADO_T64  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(CLK),
    .I(\PCI-CNTL/PCI-OFCN/PCI-XOE/NS-OE_ADO_T64 ),
    .O(OE_AD_T_T64),
    .RST(GND)
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-XOE/$5I1044  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-XOE/S_EQN64 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-XOE/B_BUSY_NS64 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/BEGIN64 )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-XOE/$5I1043  (
    .I0(B_BUSY_INT),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-XOE/$5N1033 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/B_BUSY_NS64 )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-XOE/$5I1042  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-XOE/EQN-D64 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-XOE/BH64_012 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/S_EQN64 )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-XOE/$5I1041  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$5I1041/I0 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-XOE/$5N1020 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/EQN-D64 )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-XOE/$5I1040  (
    .I0(NlwRenamedSig_OI_S_WRDN),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-XOE/$5N1019 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/END64 )
  );
  X_OR3   \PCI-CNTL/PCI-OFCN/PCI-XOE/$5I1039  (
    .I0(BH64_2),
    .I1(BH64_1),
    .I2(BH64_0),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/BH64_012 )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-XOE/$5I1038  (
    .I0(S_READY),
    .I1(S_TERM),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/$5N1020 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-OFCN/PCI-XOE/$5I1037  (
    .CE(VCC),
    .CLK(CLK),
    .I(\PCI-CNTL/PCI-OFCN/PCI-XOE/$5N1023 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/TRSTOPQ64 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-XOE/$5I1036  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-XOE/TRSTOPQ64 ),
    .I1(\FRAME- ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/$5N1019 )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-XOE/$5I1035  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$5I1035/I0 ),
    .I1(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$5I1035/I1 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/$5N1023 )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-XOE/$5I1034  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$5I1034/I0 ),
    .I1(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$5I1034/I1 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/$5N1033 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-CNTL/PCI-OFCN/PCI-XOE/OE_ADO_B  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(CLK),
    .I(\PCI-CNTL/PCI-OFCN/PCI-XOE/NS-OE_ADO_B ),
    .O(OE_AD_T_B),
    .RST(GND)
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-CNTL/PCI-OFCN/PCI-XOE/OE_ADO_T  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(CLK),
    .I(\PCI-CNTL/PCI-OFCN/PCI-XOE/NS-OE_ADO_T ),
    .O(OE_AD_T_T),
    .RST(GND)
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-CNTL/PCI-OFCN/PCI-XOE/OE_ADO_LB  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(CLK),
    .I(\PCI-CNTL/PCI-OFCN/PCI-XOE/NS-OE_ADO_LB ),
    .O(OE_AD_T_LB),
    .RST(GND)
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-CNTL/PCI-OFCN/PCI-XOE/OE_ADO_LT  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(CLK),
    .I(\PCI-CNTL/PCI-OFCN/PCI-XOE/NS-OE_ADO_LT ),
    .O(OE_AD_T_LT),
    .RST(GND)
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-XOE/$4I910  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-XOE/SET_LB ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-XOE/END ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/NS-OE_ADO_LB )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-XOE/$4I909  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$4I909/I0 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-XOE/BEGIN ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$4I909/O )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-XOE/$4I908  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$4I908/I0 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-XOE/BEGIN ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$4I908/O )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-XOE/$4I907  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-XOE/SET_LT ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-XOE/END ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/NS-OE_ADO_LT )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-XOE/$4I906  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-XOE/SET_T ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-XOE/END ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/NS-OE_ADO_T )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-XOE/$4I905  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$4I905/I0 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-XOE/BEGIN ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$4I905/O )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-XOE/$4I904  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-XOE/SET_B ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-XOE/END ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/NS-OE_ADO_B )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-XOE/$4I903  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$4I903/I0 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-XOE/BEGIN ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$4I903/O )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-XOE/$3I911  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-XOE/$3N918 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-XOE/B_BUSY_NS ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/BEGIN )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-XOE/$3I909  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-XOE/$3N905 ),
    .I1(NlwRenamedSig_OI_CFG_HIT),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/C_EQN )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-XOE/$3I900  (
    .I0(C_READY),
    .I1(C_TERM),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/$3N903 )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-XOE/$3I899  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$3I899/I0 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-XOE/$3N903 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/$3N905 )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-XOE/$3I898  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-XOE/C_EQN ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-XOE/S_EQN ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/$3N918 )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-XOE/$3I895  (
    .I0(B_BUSY_INT),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-XOE/$3N893 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/B_BUSY_NS )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-XOE/$3I890  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$3I890/I0 ),
    .I1(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$3I890/I1 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/$3N893 )
  );
  X_OR3   \PCI-CNTL/PCI-OFCN/PCI-XOE/$3I886  (
    .I0(NlwRenamedSig_OI_BASE_HIT2),
    .I1(NlwRenamedSig_OI_BASE_HIT1),
    .I2(NlwRenamedSig_OI_BASE_HIT0),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/BHIT_012 )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-XOE/$3I860  (
    .I0(NlwRenamedSig_OI_S_WRDN),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-XOE/$3N861 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/END )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CNTL/PCI-OFCN/PCI-XOE/$3I824  (
    .CE(VCC),
    .CLK(CLK),
    .I(\PCI-CNTL/PCI-OFCN/PCI-XOE/$3N818 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/TRSTOPQ ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-XOE/$3I802  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-XOE/TRSTOPQ ),
    .I1(\FRAME- ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/$3N861 )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-XOE/$3I801  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$3I801/I0 ),
    .I1(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$3I801/I1 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/$3N818 )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-XOE/$3I635  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-XOE/EQN-D ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-XOE/BHIT_012 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/S_EQN )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-XOE/$3I630  (
    .I0(S_READY),
    .I1(S_TERM),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/$3N628 )
  );
  X_OR2   \PCI-CNTL/PCI-OFCN/PCI-XOE/$3I627  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$3I627/I0 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-XOE/$3N628 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/EQN-D )
  );
  X_OR3   \PCI-CNTL/PCI-OFCN/PCI-XOE/$2I822  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-XOE/$2N1220 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-XOE/NS_HIT ),
    .I2(\PCI-CNTL/PCI-OFCN/PCI-XOE/ACTIVE ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$2I822/O )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-CNTL/PCI-OFCN/PCI-XOE/OE_DEVSEL  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(CLK),
    .I(\PCI-CNTL/PCI-OFCN/PCI-XOE/OE_TRDY_IN ),
    .O(OE_DEVSEL),
    .RST(GND)
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-CNTL/PCI-OFCN/PCI-XOE/OE_STOP  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(CLK),
    .I(\PCI-CNTL/PCI-OFCN/PCI-XOE/OE_TRDY_IN ),
    .O(OE_STOP),
    .RST(GND)
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-XOE/$2I1334  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-XOE/$2N1335 ),
    .I1(S_CYCLE64_INT),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/ACTIVE64 )
  );
  X_OR3   \PCI-CNTL/PCI-OFCN/PCI-XOE/$2I1330  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$2I1330/I0 ),
    .I1(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$2I1330/I1 ),
    .I2(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$2I1330/I2 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/$2N1335 )
  );
  X_OR3   \PCI-CNTL/PCI-OFCN/PCI-XOE/$2I1298  (
    .I0(NS_BH64_2),
    .I1(NS_BH64_1),
    .I2(NS_BH64_0),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/NS_HIT64 )
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-XOE/$2I1271  (
    .I0(B_BUSY_INT),
    .I1(\PCI-CNTL/PCI-OFCN/ACKHIT ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/$2N1272 )
  );
  X_OR3   \PCI-CNTL/PCI-OFCN/PCI-XOE/$2I1265  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-XOE/$2N1272 ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-XOE/NS_HIT64 ),
    .I2(\PCI-CNTL/PCI-OFCN/PCI-XOE/ACTIVE64 ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$2I1265/O )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-CNTL/PCI-OFCN/PCI-XOE/OE_ACK64  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(CLK),
    .I(\PCI-CNTL/PCI-OFCN/PCI-XOE/OE_ACK64_IN ),
    .O(OE_ACK64),
    .RST(GND)
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-XOE/$2I1228  (
    .I0(B_BUSY_INT),
    .I1(\PCI-CNTL/PCI-OFCN/HIT ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/$2N1220 )
  );
  X_OR4   \PCI-CNTL/PCI-OFCN/PCI-XOE/$2I1161  (
    .I0(\PCI-CNTL/NS_CFG_HIT ),
    .I1(NS_BASE_HIT2),
    .I2(NS_BASE_HIT1),
    .I3(NS_BASE_HIT0),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/NS_HIT )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-CNTL/PCI-OFCN/PCI-XOE/OE_TRDY  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(CLK),
    .I(\PCI-CNTL/PCI-OFCN/PCI-XOE/OE_TRDY_IN ),
    .O(OE_TRDY),
    .RST(GND)
  );
  X_OR3   \PCI-CNTL/PCI-OFCN/PCI-XOE/$2I1014  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$2I1014/I0 ),
    .I1(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$2I1014/I1 ),
    .I2(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$2I1014/I2 ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/ACTIVE )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-CNTL/PCI-OFCN/PCI-XOE/$1I1288  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(CLK),
    .I(\TTRDY_I- ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/TRDYDEL ),
    .RST(GND)
  );
  X_AND2   \PCI-CNTL/PCI-OFCN/PCI-XOE/$1I1270  (
    .I0(\PCI-CNTL/PCI-OFCN/PCI-XOE/HOLD_OE_PERR ),
    .I1(\PCI-CNTL/PCI-OFCN/PCI-XOE/SET_OE_PERR ),
    .O(NS_OE_PERR_T)
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-CNTL/PCI-OFCN/PCI-XOE/T_PERR_HOLD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(CLK),
    .I(\PCI-CNTL/PCI-OFCN/PCI-XOE/SET_OE_PERR ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/HOLD_OE_PERR ),
    .RST(GND)
  );
  X_AND3   \PCI-CNTL/PCI-OFCN/PCI-XOE/$1I1251  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$1I1251/I0 ),
    .I1(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$1I1251/I1 ),
    .I2(\PCI-CNTL/PCI-OFCN/PCI-XOE/EQN-A ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$1I1251/O )
  );
  X_AND4   \PCI-CNTL/PCI-OFCN/PCI-XOE/$1I1247  (
    .I0(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$1I1247/I0 ),
    .I1(NlwRenamedSig_OI_S_WRDN),
    .I2(PERR_EN),
    .I3(S_DATA_INT),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/EQN-A )
  );
  X_BUF   \PCI-CNTL/PCI-OFCN/PCI-XOE/$1I1031/NC  (
    .I(BACKOFF_INT),
    .O(\NLW_PCI-CNTL/PCI-OFCN/PCI-XOE/$1I1031/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-CNTL/PCI-OFCN/PCI-XOE/$1I1065/NC  (
    .I(TURN_AR_INT),
    .O(\NLW_PCI-CNTL/PCI-OFCN/PCI-XOE/$1I1065/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-CNTL/PCI-OFCN/PCI-XOE/$1I1239/NC  (
    .I(S_DATA_INT),
    .O(\NLW_PCI-CNTL/PCI-OFCN/PCI-XOE/$1I1239/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-CNTL/PCI-OFCN/PCI-XOE/$1I1240/NC  (
    .I(B_BUSY_INT),
    .O(\NLW_PCI-CNTL/PCI-OFCN/PCI-XOE/$1I1240/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-CNTL/$3I992/NC  (
    .I(\PCI-CNTL/TACK64- ),
    .O(\NLW_PCI-CNTL/$3I992/NC_O_UNCONNECTED )
  );
  X_AND2   \PCI-CNTL/$4I614/$1I9  (
    .I0(S_CYCLE64_INT),
    .I1(\PCI-CNTL/HOLDCYC ),
    .O(\PCI-CNTL/$4I614/M1 )
  );
  X_OR2   \PCI-CNTL/$4I614/$1I8  (
    .I0(\PCI-CNTL/$4I614/M1 ),
    .I1(\PCI-CNTL/$4I614/M0 ),
    .O(\PCI-CNTL/NS_CYC64 )
  );
  X_AND2   \PCI-CNTL/$4I614/$1I7  (
    .I0(\NlwInverterSignal_PCI-CNTL/$4I614/$1I7/I0 ),
    .I1(\PCI-CNTL/$4N752 ),
    .O(\PCI-CNTL/$4I614/M0 )
  );
  X_BUF   \$1I3754/NC  (
    .I(NlwRenamedSig_OI_ADDR31),
    .O(\NLW_$1I3754/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3755/NC  (
    .I(NlwRenamedSig_OI_ADDR30),
    .O(\NLW_$1I3755/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3756/NC  (
    .I(NlwRenamedSig_OI_ADDR29),
    .O(\NLW_$1I3756/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3757/NC  (
    .I(NlwRenamedSig_OI_ADDR28),
    .O(\NLW_$1I3757/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3758/NC  (
    .I(NlwRenamedSig_OI_ADDR27),
    .O(\NLW_$1I3758/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3759/NC  (
    .I(NlwRenamedSig_OI_ADDR26),
    .O(\NLW_$1I3759/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3760/NC  (
    .I(NlwRenamedSig_OI_ADDR25),
    .O(\NLW_$1I3760/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3761/NC  (
    .I(NlwRenamedSig_OI_ADDR24),
    .O(\NLW_$1I3761/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3762/NC  (
    .I(NlwRenamedSig_OI_ADDR23),
    .O(\NLW_$1I3762/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3763/NC  (
    .I(NlwRenamedSig_OI_ADDR22),
    .O(\NLW_$1I3763/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3764/NC  (
    .I(NlwRenamedSig_OI_ADDR21),
    .O(\NLW_$1I3764/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3765/NC  (
    .I(NlwRenamedSig_OI_ADDR20),
    .O(\NLW_$1I3765/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3766/NC  (
    .I(NlwRenamedSig_OI_ADDR19),
    .O(\NLW_$1I3766/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3767/NC  (
    .I(NlwRenamedSig_OI_ADDR18),
    .O(\NLW_$1I3767/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3768/NC  (
    .I(NlwRenamedSig_OI_ADDR17),
    .O(\NLW_$1I3768/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3769/NC  (
    .I(NlwRenamedSig_OI_ADDR16),
    .O(\NLW_$1I3769/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3770/NC  (
    .I(NlwRenamedSig_OI_ADDR15),
    .O(\NLW_$1I3770/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3771/NC  (
    .I(NlwRenamedSig_OI_ADDR14),
    .O(\NLW_$1I3771/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3772/NC  (
    .I(NlwRenamedSig_OI_ADDR13),
    .O(\NLW_$1I3772/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3773/NC  (
    .I(NlwRenamedSig_OI_ADDR12),
    .O(\NLW_$1I3773/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3774/NC  (
    .I(NlwRenamedSig_OI_ADDR11),
    .O(\NLW_$1I3774/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3775/NC  (
    .I(NlwRenamedSig_OI_ADDR10),
    .O(\NLW_$1I3775/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3776/NC  (
    .I(NlwRenamedSig_OI_ADDR9),
    .O(\NLW_$1I3776/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3777/NC  (
    .I(NlwRenamedSig_OI_ADDR8),
    .O(\NLW_$1I3777/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3778/NC  (
    .I(NlwRenamedSig_OI_ADDR7),
    .O(\NLW_$1I3778/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3779/NC  (
    .I(NlwRenamedSig_OI_ADDR6),
    .O(\NLW_$1I3779/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3780/NC  (
    .I(NlwRenamedSig_OI_ADDR5),
    .O(\NLW_$1I3780/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3781/NC  (
    .I(NlwRenamedSig_OI_ADDR4),
    .O(\NLW_$1I3781/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3782/NC  (
    .I(NlwRenamedSig_OI_ADDR3),
    .O(\NLW_$1I3782/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3783/NC  (
    .I(NlwRenamedSig_OI_ADDR2),
    .O(\NLW_$1I3783/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3784/NC  (
    .I(NlwRenamedSig_OI_ADDR1),
    .O(\NLW_$1I3784/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3785/NC  (
    .I(NlwRenamedSig_OI_ADDR0),
    .O(\NLW_$1I3785/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3786/NC  (
    .I(CE15_3),
    .O(\NLW_$1I3786/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3787/NC  (
    .I(CE15_2),
    .O(\NLW_$1I3787/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3788/NC  (
    .I(CE15_1),
    .O(\NLW_$1I3788/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3789/NC  (
    .I(CE15_0),
    .O(\NLW_$1I3789/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3790/NC  (
    .I(CE14_3),
    .O(\NLW_$1I3790/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3791/NC  (
    .I(CE14_2),
    .O(\NLW_$1I3791/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3792/NC  (
    .I(CE14_1),
    .O(\NLW_$1I3792/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3793/NC  (
    .I(CE14_0),
    .O(\NLW_$1I3793/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3794/NC  (
    .I(CE13_3),
    .O(\NLW_$1I3794/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3795/NC  (
    .I(CE13_2),
    .O(\NLW_$1I3795/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3796/NC  (
    .I(CE13_1),
    .O(\NLW_$1I3796/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3797/NC  (
    .I(CE13_0),
    .O(\NLW_$1I3797/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3798/NC  (
    .I(CE12_3),
    .O(\NLW_$1I3798/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3799/NC  (
    .I(CE12_2),
    .O(\NLW_$1I3799/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3800/NC  (
    .I(CE12_1),
    .O(\NLW_$1I3800/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3801/NC  (
    .I(CE12_0),
    .O(\NLW_$1I3801/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3802/NC  (
    .I(CE11_3),
    .O(\NLW_$1I3802/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3803/NC  (
    .I(CE11_2),
    .O(\NLW_$1I3803/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3804/NC  (
    .I(CE11_1),
    .O(\NLW_$1I3804/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3805/NC  (
    .I(CE11_0),
    .O(\NLW_$1I3805/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3806/NC  (
    .I(CE10_3),
    .O(\NLW_$1I3806/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3807/NC  (
    .I(CE10_2),
    .O(\NLW_$1I3807/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3808/NC  (
    .I(CE10_1),
    .O(\NLW_$1I3808/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3809/NC  (
    .I(CE10_0),
    .O(\NLW_$1I3809/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3810/NC  (
    .I(CE9_3),
    .O(\NLW_$1I3810/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3811/NC  (
    .I(CE9_2),
    .O(\NLW_$1I3811/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3812/NC  (
    .I(CE9_1),
    .O(\NLW_$1I3812/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3813/NC  (
    .I(CE9_0),
    .O(\NLW_$1I3813/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3814/NC  (
    .I(CE8_3),
    .O(\NLW_$1I3814/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3815/NC  (
    .I(CE8_2),
    .O(\NLW_$1I3815/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3816/NC  (
    .I(CE8_1),
    .O(\NLW_$1I3816/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3817/NC  (
    .I(CE8_0),
    .O(\NLW_$1I3817/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3818/NC  (
    .I(CE7_3),
    .O(\NLW_$1I3818/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3819/NC  (
    .I(CE7_2),
    .O(\NLW_$1I3819/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3820/NC  (
    .I(CE7_1),
    .O(\NLW_$1I3820/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3821/NC  (
    .I(CE7_0),
    .O(\NLW_$1I3821/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3822/NC  (
    .I(CE6_3),
    .O(\NLW_$1I3822/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3823/NC  (
    .I(CE6_2),
    .O(\NLW_$1I3823/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3824/NC  (
    .I(CE6_1),
    .O(\NLW_$1I3824/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3825/NC  (
    .I(CE6_0),
    .O(\NLW_$1I3825/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3826/NC  (
    .I(CE0_3),
    .O(\NLW_$1I3826/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3827/NC  (
    .I(CE0_2),
    .O(\NLW_$1I3827/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3828/NC  (
    .I(CE0_1),
    .O(\NLW_$1I3828/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3829/NC  (
    .I(CE0_0),
    .O(\NLW_$1I3829/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3830/NC  (
    .I(CE3_3),
    .O(\NLW_$1I3830/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3831/NC  (
    .I(CE3_2),
    .O(\NLW_$1I3831/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3832/NC  (
    .I(CE3_1),
    .O(\NLW_$1I3832/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3833/NC  (
    .I(CE3_0),
    .O(\NLW_$1I3833/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3834/NC  (
    .I(CE2_3),
    .O(\NLW_$1I3834/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3835/NC  (
    .I(CE2_2),
    .O(\NLW_$1I3835/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3836/NC  (
    .I(CE2_1),
    .O(\NLW_$1I3836/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3837/NC  (
    .I(CE2_0),
    .O(\NLW_$1I3837/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3840/NC  (
    .I(NlwRenamedSig_OI_PCI_CMD15),
    .O(\NLW_$1I3840/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3841/NC  (
    .I(NlwRenamedSig_OI_PCI_CMD14),
    .O(\NLW_$1I3841/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3842/NC  (
    .I(NlwRenamedSig_OI_PCI_CMD13),
    .O(\NLW_$1I3842/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3843/NC  (
    .I(NlwRenamedSig_OI_PCI_CMD12),
    .O(\NLW_$1I3843/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3844/NC  (
    .I(NlwRenamedSig_OI_PCI_CMD11),
    .O(\NLW_$1I3844/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3845/NC  (
    .I(NlwRenamedSig_OI_PCI_CMD10),
    .O(\NLW_$1I3845/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3846/NC  (
    .I(NlwRenamedSig_OI_PCI_CMD9),
    .O(\NLW_$1I3846/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3847/NC  (
    .I(NlwRenamedSig_OI_PCI_CMD8),
    .O(\NLW_$1I3847/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3848/NC  (
    .I(NlwRenamedSig_OI_PCI_CMD7),
    .O(\NLW_$1I3848/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3849/NC  (
    .I(NlwRenamedSig_OI_PCI_CMD6),
    .O(\NLW_$1I3849/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3850/NC  (
    .I(NlwRenamedSig_OI_PCI_CMD5),
    .O(\NLW_$1I3850/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3851/NC  (
    .I(NlwRenamedSig_OI_PCI_CMD4),
    .O(\NLW_$1I3851/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3852/NC  (
    .I(NlwRenamedSig_OI_PCI_CMD3),
    .O(\NLW_$1I3852/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3853/NC  (
    .I(NlwRenamedSig_OI_PCI_CMD2),
    .O(\NLW_$1I3853/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3854/NC  (
    .I(NlwRenamedSig_OI_PCI_CMD1),
    .O(\NLW_$1I3854/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3855/NC  (
    .I(NlwRenamedSig_OI_PCI_CMD0),
    .O(\NLW_$1I3855/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3860/NC  (
    .I(OE15),
    .O(\NLW_$1I3860/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3861/NC  (
    .I(OE14),
    .O(\NLW_$1I3861/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3862/NC  (
    .I(OE13),
    .O(\NLW_$1I3862/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3863/NC  (
    .I(OE12),
    .O(\NLW_$1I3863/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3864/NC  (
    .I(OE11),
    .O(\NLW_$1I3864/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3865/NC  (
    .I(OE10),
    .O(\NLW_$1I3865/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3866/NC  (
    .I(OE9),
    .O(\NLW_$1I3866/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3867/NC  (
    .I(OE8),
    .O(\NLW_$1I3867/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3868/NC  (
    .I(OE7),
    .O(\NLW_$1I3868/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3869/NC  (
    .I(OE6),
    .O(\NLW_$1I3869/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3870/NC  (
    .I(OE5),
    .O(\NLW_$1I3870/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3871/NC  (
    .I(OE4),
    .O(\NLW_$1I3871/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3872/NC  (
    .I(OE3),
    .O(\NLW_$1I3872/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3873/NC  (
    .I(OE2),
    .O(\NLW_$1I3873/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3874/NC  (
    .I(OE1),
    .O(\NLW_$1I3874/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3875/NC  (
    .I(OE0),
    .O(\NLW_$1I3875/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3879/NC  (
    .I(NlwRenamedSig_OI_CSR39),
    .O(\NLW_$1I3879/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3880/NC  (
    .I(NlwRenamedSig_OI_CSR38),
    .O(\NLW_$1I3880/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3881/NC  (
    .I(NlwRenamedSig_OI_CSR37),
    .O(\NLW_$1I3881/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3882/NC  (
    .I(NlwRenamedSig_OI_CSR36),
    .O(\NLW_$1I3882/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3883/NC  (
    .I(NlwRenamedSig_OI_CSR35),
    .O(\NLW_$1I3883/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3884/NC  (
    .I(NlwRenamedSig_OI_CSR34),
    .O(\NLW_$1I3884/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3885/NC  (
    .I(NlwRenamedSig_OI_CSR33),
    .O(\NLW_$1I3885/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3886/NC  (
    .I(NlwRenamedSig_OI_CSR32),
    .O(\NLW_$1I3886/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3887/NC  (
    .I(NlwRenamedSig_OI_CSR31),
    .O(\NLW_$1I3887/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3888/NC  (
    .I(NlwRenamedSig_OI_CSR30),
    .O(\NLW_$1I3888/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3889/NC  (
    .I(NlwRenamedSig_OI_CSR29),
    .O(\NLW_$1I3889/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3890/NC  (
    .I(NlwRenamedSig_OI_CSR28),
    .O(\NLW_$1I3890/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3891/NC  (
    .I(NlwRenamedSig_OI_CSR27),
    .O(\NLW_$1I3891/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3892/NC  (
    .I(NlwRenamedSig_OI_CSR26),
    .O(\NLW_$1I3892/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3893/NC  (
    .I(NlwRenamedSig_OI_CSR25),
    .O(\NLW_$1I3893/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3894/NC  (
    .I(NlwRenamedSig_OI_CSR24),
    .O(\NLW_$1I3894/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3895/NC  (
    .I(NlwRenamedSig_OI_CSR23),
    .O(\NLW_$1I3895/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3896/NC  (
    .I(NlwRenamedSig_OI_CSR22),
    .O(\NLW_$1I3896/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3897/NC  (
    .I(NlwRenamedSig_OI_CSR21),
    .O(\NLW_$1I3897/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3898/NC  (
    .I(NlwRenamedSig_OI_CSR20),
    .O(\NLW_$1I3898/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3899/NC  (
    .I(NlwRenamedSig_OI_CSR19),
    .O(\NLW_$1I3899/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3900/NC  (
    .I(NlwRenamedSig_OI_CSR18),
    .O(\NLW_$1I3900/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3901/NC  (
    .I(NlwRenamedSig_OI_CSR17),
    .O(\NLW_$1I3901/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3902/NC  (
    .I(NlwRenamedSig_OI_CSR16),
    .O(\NLW_$1I3902/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3903/NC  (
    .I(NlwRenamedSig_OI_CSR15),
    .O(\NLW_$1I3903/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3904/NC  (
    .I(NlwRenamedSig_OI_CSR14),
    .O(\NLW_$1I3904/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3905/NC  (
    .I(NlwRenamedSig_OI_CSR13),
    .O(\NLW_$1I3905/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3906/NC  (
    .I(NlwRenamedSig_OI_CSR12),
    .O(\NLW_$1I3906/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3907/NC  (
    .I(NlwRenamedSig_OI_CSR11),
    .O(\NLW_$1I3907/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3908/NC  (
    .I(NlwRenamedSig_OI_CSR10),
    .O(\NLW_$1I3908/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3909/NC  (
    .I(NlwRenamedSig_OI_CSR9),
    .O(\NLW_$1I3909/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3910/NC  (
    .I(NlwRenamedSig_OI_CSR8),
    .O(\NLW_$1I3910/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3911/NC  (
    .I(NlwRenamedSig_OI_CSR7),
    .O(\NLW_$1I3911/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3912/NC  (
    .I(NlwRenamedSig_OI_CSR6),
    .O(\NLW_$1I3912/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3913/NC  (
    .I(NlwRenamedSig_OI_CSR5),
    .O(\NLW_$1I3913/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3914/NC  (
    .I(NlwRenamedSig_OI_CSR4),
    .O(\NLW_$1I3914/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3915/NC  (
    .I(NlwRenamedSig_OI_CSR3),
    .O(\NLW_$1I3915/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3916/NC  (
    .I(NlwRenamedSig_OI_CSR2),
    .O(\NLW_$1I3916/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3917/NC  (
    .I(NlwRenamedSig_OI_CSR1),
    .O(\NLW_$1I3917/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3918/NC  (
    .I(NlwRenamedSig_OI_CSR0),
    .O(\NLW_$1I3918/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3921/NC  (
    .I(NlwRenamedSig_OI_S_CBE7),
    .O(\NLW_$1I3921/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3922/NC  (
    .I(NlwRenamedSig_OI_S_CBE6),
    .O(\NLW_$1I3922/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3923/NC  (
    .I(NlwRenamedSig_OI_S_CBE5),
    .O(\NLW_$1I3923/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3924/NC  (
    .I(NlwRenamedSig_OI_S_CBE4),
    .O(\NLW_$1I3924/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3925/NC  (
    .I(NlwRenamedSig_OI_S_CBE3),
    .O(\NLW_$1I3925/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3926/NC  (
    .I(NlwRenamedSig_OI_S_CBE2),
    .O(\NLW_$1I3926/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3927/NC  (
    .I(NlwRenamedSig_OI_S_CBE1),
    .O(\NLW_$1I3927/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I3928/NC  (
    .I(NlwRenamedSig_OI_S_CBE0),
    .O(\NLW_$1I3928/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4355/NC  (
    .I(CFG255),
    .O(\NLW_$1I4355/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4356/NC  (
    .I(CFG254),
    .O(\NLW_$1I4356/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4357/NC  (
    .I(CFG253),
    .O(\NLW_$1I4357/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4358/NC  (
    .I(CFG252),
    .O(\NLW_$1I4358/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4359/NC  (
    .I(CFG251),
    .O(\NLW_$1I4359/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4360/NC  (
    .I(CFG250),
    .O(\NLW_$1I4360/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4361/NC  (
    .I(CFG249),
    .O(\NLW_$1I4361/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4362/NC  (
    .I(CFG248),
    .O(\NLW_$1I4362/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4363/NC  (
    .I(CFG247),
    .O(\NLW_$1I4363/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4364/NC  (
    .I(CFG246),
    .O(\NLW_$1I4364/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4365/NC  (
    .I(CFG245),
    .O(\NLW_$1I4365/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4366/NC  (
    .I(CFG244),
    .O(\NLW_$1I4366/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4367/NC  (
    .I(CFG243),
    .O(\NLW_$1I4367/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4368/NC  (
    .I(CFG242),
    .O(\NLW_$1I4368/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4369/NC  (
    .I(CFG241),
    .O(\NLW_$1I4369/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4370/NC  (
    .I(CFG240),
    .O(\NLW_$1I4370/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4371/NC  (
    .I(CFG239),
    .O(\NLW_$1I4371/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4372/NC  (
    .I(CFG238),
    .O(\NLW_$1I4372/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4373/NC  (
    .I(CFG237),
    .O(\NLW_$1I4373/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4374/NC  (
    .I(CFG236),
    .O(\NLW_$1I4374/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4375/NC  (
    .I(CFG235),
    .O(\NLW_$1I4375/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4376/NC  (
    .I(CFG234),
    .O(\NLW_$1I4376/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4377/NC  (
    .I(CFG233),
    .O(\NLW_$1I4377/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4378/NC  (
    .I(CFG232),
    .O(\NLW_$1I4378/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4379/NC  (
    .I(CFG231),
    .O(\NLW_$1I4379/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4380/NC  (
    .I(CFG230),
    .O(\NLW_$1I4380/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4381/NC  (
    .I(CFG229),
    .O(\NLW_$1I4381/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4382/NC  (
    .I(CFG228),
    .O(\NLW_$1I4382/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4383/NC  (
    .I(CFG227),
    .O(\NLW_$1I4383/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4384/NC  (
    .I(CFG226),
    .O(\NLW_$1I4384/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4385/NC  (
    .I(CFG225),
    .O(\NLW_$1I4385/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4386/NC  (
    .I(CFG224),
    .O(\NLW_$1I4386/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4387/NC  (
    .I(CFG223),
    .O(\NLW_$1I4387/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4388/NC  (
    .I(CFG222),
    .O(\NLW_$1I4388/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4389/NC  (
    .I(CFG221),
    .O(\NLW_$1I4389/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4390/NC  (
    .I(CFG220),
    .O(\NLW_$1I4390/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4391/NC  (
    .I(CFG219),
    .O(\NLW_$1I4391/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4392/NC  (
    .I(CFG218),
    .O(\NLW_$1I4392/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4393/NC  (
    .I(CFG217),
    .O(\NLW_$1I4393/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4394/NC  (
    .I(CFG216),
    .O(\NLW_$1I4394/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4395/NC  (
    .I(CFG215),
    .O(\NLW_$1I4395/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4396/NC  (
    .I(CFG214),
    .O(\NLW_$1I4396/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4397/NC  (
    .I(CFG213),
    .O(\NLW_$1I4397/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4398/NC  (
    .I(CFG212),
    .O(\NLW_$1I4398/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4399/NC  (
    .I(CFG211),
    .O(\NLW_$1I4399/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4400/NC  (
    .I(CFG210),
    .O(\NLW_$1I4400/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4401/NC  (
    .I(CFG209),
    .O(\NLW_$1I4401/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4402/NC  (
    .I(CFG208),
    .O(\NLW_$1I4402/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4403/NC  (
    .I(CFG207),
    .O(\NLW_$1I4403/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4404/NC  (
    .I(CFG206),
    .O(\NLW_$1I4404/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4405/NC  (
    .I(CFG205),
    .O(\NLW_$1I4405/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4406/NC  (
    .I(CFG204),
    .O(\NLW_$1I4406/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4407/NC  (
    .I(CFG203),
    .O(\NLW_$1I4407/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4408/NC  (
    .I(CFG202),
    .O(\NLW_$1I4408/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4409/NC  (
    .I(CFG201),
    .O(\NLW_$1I4409/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4410/NC  (
    .I(CFG200),
    .O(\NLW_$1I4410/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4411/NC  (
    .I(CFG199),
    .O(\NLW_$1I4411/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4412/NC  (
    .I(CFG198),
    .O(\NLW_$1I4412/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4413/NC  (
    .I(CFG197),
    .O(\NLW_$1I4413/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4414/NC  (
    .I(CFG196),
    .O(\NLW_$1I4414/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4415/NC  (
    .I(CFG195),
    .O(\NLW_$1I4415/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4416/NC  (
    .I(CFG194),
    .O(\NLW_$1I4416/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4417/NC  (
    .I(CFG193),
    .O(\NLW_$1I4417/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4418/NC  (
    .I(CFG192),
    .O(\NLW_$1I4418/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4419/NC  (
    .I(CFG191),
    .O(\NLW_$1I4419/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4420/NC  (
    .I(CFG190),
    .O(\NLW_$1I4420/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4421/NC  (
    .I(CFG189),
    .O(\NLW_$1I4421/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4422/NC  (
    .I(CFG188),
    .O(\NLW_$1I4422/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4423/NC  (
    .I(CFG187),
    .O(\NLW_$1I4423/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4424/NC  (
    .I(CFG186),
    .O(\NLW_$1I4424/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4425/NC  (
    .I(CFG185),
    .O(\NLW_$1I4425/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4426/NC  (
    .I(CFG184),
    .O(\NLW_$1I4426/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4427/NC  (
    .I(CFG183),
    .O(\NLW_$1I4427/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4428/NC  (
    .I(CFG182),
    .O(\NLW_$1I4428/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4429/NC  (
    .I(CFG181),
    .O(\NLW_$1I4429/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4430/NC  (
    .I(CFG180),
    .O(\NLW_$1I4430/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4431/NC  (
    .I(CFG179),
    .O(\NLW_$1I4431/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4432/NC  (
    .I(CFG178),
    .O(\NLW_$1I4432/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4433/NC  (
    .I(CFG177),
    .O(\NLW_$1I4433/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4434/NC  (
    .I(CFG176),
    .O(\NLW_$1I4434/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4435/NC  (
    .I(CFG175),
    .O(\NLW_$1I4435/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4436/NC  (
    .I(CFG174),
    .O(\NLW_$1I4436/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4437/NC  (
    .I(CFG173),
    .O(\NLW_$1I4437/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4438/NC  (
    .I(CFG172),
    .O(\NLW_$1I4438/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4439/NC  (
    .I(CFG171),
    .O(\NLW_$1I4439/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4440/NC  (
    .I(CFG170),
    .O(\NLW_$1I4440/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4441/NC  (
    .I(CFG169),
    .O(\NLW_$1I4441/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4442/NC  (
    .I(CFG168),
    .O(\NLW_$1I4442/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4443/NC  (
    .I(CFG167),
    .O(\NLW_$1I4443/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4444/NC  (
    .I(CFG166),
    .O(\NLW_$1I4444/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4445/NC  (
    .I(CFG165),
    .O(\NLW_$1I4445/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4446/NC  (
    .I(CFG164),
    .O(\NLW_$1I4446/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4447/NC  (
    .I(CFG163),
    .O(\NLW_$1I4447/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4448/NC  (
    .I(CFG162),
    .O(\NLW_$1I4448/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4449/NC  (
    .I(CFG161),
    .O(\NLW_$1I4449/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4450/NC  (
    .I(CFG160),
    .O(\NLW_$1I4450/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4451/NC  (
    .I(CFG159),
    .O(\NLW_$1I4451/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4452/NC  (
    .I(CFG158),
    .O(\NLW_$1I4452/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4453/NC  (
    .I(CFG157),
    .O(\NLW_$1I4453/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4454/NC  (
    .I(CFG156),
    .O(\NLW_$1I4454/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4455/NC  (
    .I(CFG155),
    .O(\NLW_$1I4455/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4456/NC  (
    .I(CFG154),
    .O(\NLW_$1I4456/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4457/NC  (
    .I(CFG153),
    .O(\NLW_$1I4457/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4458/NC  (
    .I(CFG152),
    .O(\NLW_$1I4458/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4459/NC  (
    .I(CFG151),
    .O(\NLW_$1I4459/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4460/NC  (
    .I(CFG150),
    .O(\NLW_$1I4460/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4461/NC  (
    .I(CFG149),
    .O(\NLW_$1I4461/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4462/NC  (
    .I(CFG148),
    .O(\NLW_$1I4462/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4463/NC  (
    .I(CFG147),
    .O(\NLW_$1I4463/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4464/NC  (
    .I(CFG146),
    .O(\NLW_$1I4464/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4465/NC  (
    .I(CFG145),
    .O(\NLW_$1I4465/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4466/NC  (
    .I(CFG144),
    .O(\NLW_$1I4466/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4467/NC  (
    .I(CFG143),
    .O(\NLW_$1I4467/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4468/NC  (
    .I(CFG142),
    .O(\NLW_$1I4468/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4469/NC  (
    .I(CFG141),
    .O(\NLW_$1I4469/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4470/NC  (
    .I(CFG140),
    .O(\NLW_$1I4470/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4471/NC  (
    .I(CFG139),
    .O(\NLW_$1I4471/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4472/NC  (
    .I(CFG138),
    .O(\NLW_$1I4472/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4473/NC  (
    .I(CFG137),
    .O(\NLW_$1I4473/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4474/NC  (
    .I(CFG136),
    .O(\NLW_$1I4474/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4475/NC  (
    .I(CFG135),
    .O(\NLW_$1I4475/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4476/NC  (
    .I(CFG134),
    .O(\NLW_$1I4476/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4477/NC  (
    .I(CFG133),
    .O(\NLW_$1I4477/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4478/NC  (
    .I(CFG132),
    .O(\NLW_$1I4478/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4479/NC  (
    .I(CFG131),
    .O(\NLW_$1I4479/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4480/NC  (
    .I(CFG130),
    .O(\NLW_$1I4480/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4481/NC  (
    .I(CFG129),
    .O(\NLW_$1I4481/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4482/NC  (
    .I(CFG128),
    .O(\NLW_$1I4482/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4483/NC  (
    .I(CFG127),
    .O(\NLW_$1I4483/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4484/NC  (
    .I(CFG126),
    .O(\NLW_$1I4484/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4485/NC  (
    .I(CFG125),
    .O(\NLW_$1I4485/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4486/NC  (
    .I(CFG124),
    .O(\NLW_$1I4486/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4487/NC  (
    .I(CFG123),
    .O(\NLW_$1I4487/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4488/NC  (
    .I(CFG122),
    .O(\NLW_$1I4488/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4489/NC  (
    .I(CFG121),
    .O(\NLW_$1I4489/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4490/NC  (
    .I(CFG120),
    .O(\NLW_$1I4490/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4491/NC  (
    .I(CFG119),
    .O(\NLW_$1I4491/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4492/NC  (
    .I(CFG118),
    .O(\NLW_$1I4492/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4493/NC  (
    .I(CFG117),
    .O(\NLW_$1I4493/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4494/NC  (
    .I(CFG116),
    .O(\NLW_$1I4494/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4495/NC  (
    .I(CFG115),
    .O(\NLW_$1I4495/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4496/NC  (
    .I(CFG114),
    .O(\NLW_$1I4496/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4497/NC  (
    .I(CFG113),
    .O(\NLW_$1I4497/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4498/NC  (
    .I(CFG112),
    .O(\NLW_$1I4498/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4499/NC  (
    .I(CFG111),
    .O(\NLW_$1I4499/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4500/NC  (
    .I(CFG110),
    .O(\NLW_$1I4500/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4501/NC  (
    .I(CFG109),
    .O(\NLW_$1I4501/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4502/NC  (
    .I(CFG108),
    .O(\NLW_$1I4502/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4503/NC  (
    .I(CFG107),
    .O(\NLW_$1I4503/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4504/NC  (
    .I(CFG106),
    .O(\NLW_$1I4504/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4505/NC  (
    .I(CFG105),
    .O(\NLW_$1I4505/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4506/NC  (
    .I(CFG104),
    .O(\NLW_$1I4506/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4507/NC  (
    .I(CFG103),
    .O(\NLW_$1I4507/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4508/NC  (
    .I(CFG102),
    .O(\NLW_$1I4508/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4509/NC  (
    .I(CFG101),
    .O(\NLW_$1I4509/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4510/NC  (
    .I(CFG100),
    .O(\NLW_$1I4510/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4511/NC  (
    .I(CFG99),
    .O(\NLW_$1I4511/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4512/NC  (
    .I(CFG98),
    .O(\NLW_$1I4512/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4513/NC  (
    .I(CFG97),
    .O(\NLW_$1I4513/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4514/NC  (
    .I(CFG96),
    .O(\NLW_$1I4514/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4515/NC  (
    .I(CFG95),
    .O(\NLW_$1I4515/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4516/NC  (
    .I(CFG94),
    .O(\NLW_$1I4516/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4517/NC  (
    .I(CFG93),
    .O(\NLW_$1I4517/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4518/NC  (
    .I(CFG92),
    .O(\NLW_$1I4518/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4519/NC  (
    .I(CFG91),
    .O(\NLW_$1I4519/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4520/NC  (
    .I(CFG90),
    .O(\NLW_$1I4520/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4521/NC  (
    .I(CFG89),
    .O(\NLW_$1I4521/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4522/NC  (
    .I(CFG88),
    .O(\NLW_$1I4522/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4523/NC  (
    .I(CFG87),
    .O(\NLW_$1I4523/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4524/NC  (
    .I(CFG86),
    .O(\NLW_$1I4524/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4525/NC  (
    .I(CFG85),
    .O(\NLW_$1I4525/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4526/NC  (
    .I(CFG84),
    .O(\NLW_$1I4526/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4527/NC  (
    .I(CFG83),
    .O(\NLW_$1I4527/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4528/NC  (
    .I(CFG82),
    .O(\NLW_$1I4528/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4529/NC  (
    .I(CFG81),
    .O(\NLW_$1I4529/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4530/NC  (
    .I(CFG80),
    .O(\NLW_$1I4530/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4531/NC  (
    .I(CFG79),
    .O(\NLW_$1I4531/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4532/NC  (
    .I(CFG78),
    .O(\NLW_$1I4532/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4533/NC  (
    .I(CFG77),
    .O(\NLW_$1I4533/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4534/NC  (
    .I(CFG76),
    .O(\NLW_$1I4534/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4535/NC  (
    .I(CFG75),
    .O(\NLW_$1I4535/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4536/NC  (
    .I(CFG74),
    .O(\NLW_$1I4536/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4537/NC  (
    .I(CFG73),
    .O(\NLW_$1I4537/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4538/NC  (
    .I(CFG72),
    .O(\NLW_$1I4538/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4539/NC  (
    .I(CFG71),
    .O(\NLW_$1I4539/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4540/NC  (
    .I(CFG70),
    .O(\NLW_$1I4540/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4541/NC  (
    .I(CFG69),
    .O(\NLW_$1I4541/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4542/NC  (
    .I(CFG68),
    .O(\NLW_$1I4542/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4543/NC  (
    .I(CFG67),
    .O(\NLW_$1I4543/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4544/NC  (
    .I(CFG66),
    .O(\NLW_$1I4544/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4545/NC  (
    .I(CFG65),
    .O(\NLW_$1I4545/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4546/NC  (
    .I(CFG64),
    .O(\NLW_$1I4546/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4547/NC  (
    .I(CFG63),
    .O(\NLW_$1I4547/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4548/NC  (
    .I(CFG62),
    .O(\NLW_$1I4548/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4549/NC  (
    .I(CFG61),
    .O(\NLW_$1I4549/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4550/NC  (
    .I(CFG60),
    .O(\NLW_$1I4550/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4551/NC  (
    .I(CFG59),
    .O(\NLW_$1I4551/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4552/NC  (
    .I(CFG58),
    .O(\NLW_$1I4552/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4553/NC  (
    .I(CFG57),
    .O(\NLW_$1I4553/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4554/NC  (
    .I(CFG56),
    .O(\NLW_$1I4554/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4555/NC  (
    .I(CFG55),
    .O(\NLW_$1I4555/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4556/NC  (
    .I(CFG54),
    .O(\NLW_$1I4556/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4557/NC  (
    .I(CFG53),
    .O(\NLW_$1I4557/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4558/NC  (
    .I(CFG52),
    .O(\NLW_$1I4558/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4559/NC  (
    .I(CFG51),
    .O(\NLW_$1I4559/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4560/NC  (
    .I(CFG50),
    .O(\NLW_$1I4560/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4561/NC  (
    .I(CFG49),
    .O(\NLW_$1I4561/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4562/NC  (
    .I(CFG48),
    .O(\NLW_$1I4562/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4563/NC  (
    .I(CFG47),
    .O(\NLW_$1I4563/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4564/NC  (
    .I(CFG46),
    .O(\NLW_$1I4564/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4565/NC  (
    .I(CFG45),
    .O(\NLW_$1I4565/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4566/NC  (
    .I(CFG44),
    .O(\NLW_$1I4566/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4567/NC  (
    .I(CFG43),
    .O(\NLW_$1I4567/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4568/NC  (
    .I(CFG42),
    .O(\NLW_$1I4568/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4569/NC  (
    .I(CFG41),
    .O(\NLW_$1I4569/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4570/NC  (
    .I(CFG40),
    .O(\NLW_$1I4570/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4571/NC  (
    .I(CFG39),
    .O(\NLW_$1I4571/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4572/NC  (
    .I(CFG38),
    .O(\NLW_$1I4572/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4573/NC  (
    .I(CFG37),
    .O(\NLW_$1I4573/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4574/NC  (
    .I(CFG36),
    .O(\NLW_$1I4574/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4575/NC  (
    .I(CFG35),
    .O(\NLW_$1I4575/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4576/NC  (
    .I(CFG34),
    .O(\NLW_$1I4576/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4577/NC  (
    .I(CFG33),
    .O(\NLW_$1I4577/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4578/NC  (
    .I(CFG32),
    .O(\NLW_$1I4578/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4579/NC  (
    .I(CFG31),
    .O(\NLW_$1I4579/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4580/NC  (
    .I(CFG30),
    .O(\NLW_$1I4580/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4581/NC  (
    .I(CFG29),
    .O(\NLW_$1I4581/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4582/NC  (
    .I(CFG28),
    .O(\NLW_$1I4582/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4583/NC  (
    .I(CFG27),
    .O(\NLW_$1I4583/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4584/NC  (
    .I(CFG26),
    .O(\NLW_$1I4584/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4585/NC  (
    .I(CFG25),
    .O(\NLW_$1I4585/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4586/NC  (
    .I(CFG24),
    .O(\NLW_$1I4586/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4587/NC  (
    .I(CFG23),
    .O(\NLW_$1I4587/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4588/NC  (
    .I(CFG22),
    .O(\NLW_$1I4588/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4589/NC  (
    .I(CFG21),
    .O(\NLW_$1I4589/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4590/NC  (
    .I(CFG20),
    .O(\NLW_$1I4590/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4591/NC  (
    .I(CFG19),
    .O(\NLW_$1I4591/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4592/NC  (
    .I(CFG18),
    .O(\NLW_$1I4592/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4593/NC  (
    .I(CFG17),
    .O(\NLW_$1I4593/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4594/NC  (
    .I(CFG16),
    .O(\NLW_$1I4594/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4595/NC  (
    .I(CFG15),
    .O(\NLW_$1I4595/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4596/NC  (
    .I(CFG14),
    .O(\NLW_$1I4596/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4597/NC  (
    .I(CFG13),
    .O(\NLW_$1I4597/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4598/NC  (
    .I(CFG12),
    .O(\NLW_$1I4598/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4599/NC  (
    .I(CFG11),
    .O(\NLW_$1I4599/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4600/NC  (
    .I(CFG10),
    .O(\NLW_$1I4600/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4601/NC  (
    .I(CFG9),
    .O(\NLW_$1I4601/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4602/NC  (
    .I(CFG8),
    .O(\NLW_$1I4602/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4603/NC  (
    .I(CFG7),
    .O(\NLW_$1I4603/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4604/NC  (
    .I(CFG6),
    .O(\NLW_$1I4604/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4605/NC  (
    .I(CFG5),
    .O(\NLW_$1I4605/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4606/NC  (
    .I(CFG4),
    .O(\NLW_$1I4606/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4607/NC  (
    .I(CFG3),
    .O(\NLW_$1I4607/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4608/NC  (
    .I(CFG2),
    .O(\NLW_$1I4608/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4609/NC  (
    .I(CFG1),
    .O(\NLW_$1I4609/NC_O_UNCONNECTED )
  );
  X_BUF   \$1I4610/NC  (
    .I(CFG0),
    .O(\NLW_$1I4610/NC_O_UNCONNECTED )
  );
  X_BUF   \TDLY/$1I269  (
    .I(\TDLY/D5_4117 ),
    .O(\TDLY/D6_4118 )
  );
  X_BUF   \TDLY/$1I266  (
    .I(\TDLY/D4_4116 ),
    .O(\TDLY/D5_4117 )
  );
  X_BUF   \TDLY/$1I255  (
    .I(\TDLY/D3_4115 ),
    .O(\TDLY/D4_4116 )
  );
  X_BUF   \TDLY/$1I251  (
    .I(\TDLY/D2_4114 ),
    .O(\TDLY/D3_4115 )
  );
  X_BUF   \TDLY/$1I245  (
    .I(\TDLY/D1_4113 ),
    .O(\TDLY/D2_4114 )
  );
  X_BUF   \TDLY/$1I236  (
    .I(TRDY_I),
    .O(\TDLY/D1_4113 )
  );
  X_MUX2   \TDLY/$1I315/O  (
    .IA(\TDLY/$1I315/M01 ),
    .IB(\TDLY/$1I315/M23 ),
    .O(TRDY_F),
    .SEL(CFG246)
  );
  X_OR2   \TDLY/$1I315/M01/$1I38  (
    .I0(\TDLY/$1I315/M01/M1 ),
    .I1(\TDLY/$1I315/M01/M0 ),
    .O(\TDLY/$1I315/M01 )
  );
  X_AND3   \TDLY/$1I315/M01/$1I31  (
    .I0(\NlwInverterSignal_TDLY/$1I315/M01/$1I31/I0 ),
    .I1(\TDLY/$1N318 ),
    .I2(TRDY_I),
    .O(\TDLY/$1I315/M01/M0 )
  );
  X_AND3   \TDLY/$1I315/M01/$1I30  (
    .I0(\TDLY/D1_4113 ),
    .I1(\TDLY/$1N318 ),
    .I2(CFG245),
    .O(\TDLY/$1I315/M01/M1 )
  );
  X_OR2   \TDLY/$1I315/M23/$1I38  (
    .I0(\TDLY/$1I315/M23/M1 ),
    .I1(\TDLY/$1I315/M23/M0 ),
    .O(\TDLY/$1I315/M23 )
  );
  X_AND3   \TDLY/$1I315/M23/$1I31  (
    .I0(\NlwInverterSignal_TDLY/$1I315/M23/$1I31/I0 ),
    .I1(\TDLY/$1N318 ),
    .I2(\TDLY/D2_4114 ),
    .O(\TDLY/$1I315/M23/M0 )
  );
  X_AND3   \TDLY/$1I315/M23/$1I30  (
    .I0(\TDLY/D3_4115 ),
    .I1(\TDLY/$1N318 ),
    .I2(CFG245),
    .O(\TDLY/$1I315/M23/M1 )
  );
  X_ONE   \TDLY/$1I319/$1I2220  (
    .O(\TDLY/$1I319/$1N2216 )
  );
  X_BUF   \TDLY/$1I319/H  (
    .I(\TDLY/$1I319/$1N2216 ),
    .O(\TDLY/$1N318 )
  );
  X_MUX2   \TDLY/$1I328/O  (
    .IA(\TDLY/$1I328/M01 ),
    .IB(\TDLY/$1I328/M23 ),
    .O(TRDY_M),
    .SEL(CFG246)
  );
  X_OR2   \TDLY/$1I328/M01/$1I38  (
    .I0(\TDLY/$1I328/M01/M1 ),
    .I1(\TDLY/$1I328/M01/M0 ),
    .O(\TDLY/$1I328/M01 )
  );
  X_AND3   \TDLY/$1I328/M01/$1I31  (
    .I0(\NlwInverterSignal_TDLY/$1I328/M01/$1I31/I0 ),
    .I1(\TDLY/$1N332 ),
    .I2(TRDY_I),
    .O(\TDLY/$1I328/M01/M0 )
  );
  X_AND3   \TDLY/$1I328/M01/$1I30  (
    .I0(\TDLY/D3_4115 ),
    .I1(\TDLY/$1N332 ),
    .I2(CFG245),
    .O(\TDLY/$1I328/M01/M1 )
  );
  X_OR2   \TDLY/$1I328/M23/$1I38  (
    .I0(\TDLY/$1I328/M23/M1 ),
    .I1(\TDLY/$1I328/M23/M0 ),
    .O(\TDLY/$1I328/M23 )
  );
  X_AND3   \TDLY/$1I328/M23/$1I31  (
    .I0(\NlwInverterSignal_TDLY/$1I328/M23/$1I31/I0 ),
    .I1(\TDLY/$1N332 ),
    .I2(\TDLY/D4_4116 ),
    .O(\TDLY/$1I328/M23/M0 )
  );
  X_AND3   \TDLY/$1I328/M23/$1I30  (
    .I0(\TDLY/D5_4117 ),
    .I1(\TDLY/$1N332 ),
    .I2(CFG245),
    .O(\TDLY/$1I328/M23/M1 )
  );
  X_ONE   \TDLY/$1I331/$1I2220  (
    .O(\TDLY/$1I331/$1N2216 )
  );
  X_BUF   \TDLY/$1I331/H  (
    .I(\TDLY/$1I331/$1N2216 ),
    .O(\TDLY/$1N332 )
  );
  X_BUF   \IDLY/$1I269  (
    .I(\IDLY/D5_4182 ),
    .O(\IDLY/D6_4183 )
  );
  X_BUF   \IDLY/$1I266  (
    .I(\IDLY/D4_4181 ),
    .O(\IDLY/D5_4182 )
  );
  X_BUF   \IDLY/$1I255  (
    .I(\IDLY/D3_4180 ),
    .O(\IDLY/D4_4181 )
  );
  X_BUF   \IDLY/$1I251  (
    .I(\IDLY/D2_4179 ),
    .O(\IDLY/D3_4180 )
  );
  X_BUF   \IDLY/$1I245  (
    .I(\IDLY/D1_4178 ),
    .O(\IDLY/D2_4179 )
  );
  X_BUF   \IDLY/$1I236  (
    .I(IRDY_I),
    .O(\IDLY/D1_4178 )
  );
  X_MUX2   \IDLY/$1I315/O  (
    .IA(\IDLY/$1I315/M01 ),
    .IB(\IDLY/$1I315/M23 ),
    .O(IRDY_F),
    .SEL(CFG246)
  );
  X_OR2   \IDLY/$1I315/M01/$1I38  (
    .I0(\IDLY/$1I315/M01/M1 ),
    .I1(\IDLY/$1I315/M01/M0 ),
    .O(\IDLY/$1I315/M01 )
  );
  X_AND3   \IDLY/$1I315/M01/$1I31  (
    .I0(\NlwInverterSignal_IDLY/$1I315/M01/$1I31/I0 ),
    .I1(\IDLY/$1N318 ),
    .I2(IRDY_I),
    .O(\IDLY/$1I315/M01/M0 )
  );
  X_AND3   \IDLY/$1I315/M01/$1I30  (
    .I0(\IDLY/D1_4178 ),
    .I1(\IDLY/$1N318 ),
    .I2(CFG245),
    .O(\IDLY/$1I315/M01/M1 )
  );
  X_OR2   \IDLY/$1I315/M23/$1I38  (
    .I0(\IDLY/$1I315/M23/M1 ),
    .I1(\IDLY/$1I315/M23/M0 ),
    .O(\IDLY/$1I315/M23 )
  );
  X_AND3   \IDLY/$1I315/M23/$1I31  (
    .I0(\NlwInverterSignal_IDLY/$1I315/M23/$1I31/I0 ),
    .I1(\IDLY/$1N318 ),
    .I2(\IDLY/D2_4179 ),
    .O(\IDLY/$1I315/M23/M0 )
  );
  X_AND3   \IDLY/$1I315/M23/$1I30  (
    .I0(\IDLY/D3_4180 ),
    .I1(\IDLY/$1N318 ),
    .I2(CFG245),
    .O(\IDLY/$1I315/M23/M1 )
  );
  X_ONE   \IDLY/$1I319/$1I2220  (
    .O(\IDLY/$1I319/$1N2216 )
  );
  X_BUF   \IDLY/$1I319/H  (
    .I(\IDLY/$1I319/$1N2216 ),
    .O(\IDLY/$1N318 )
  );
  X_MUX2   \IDLY/$1I328/O  (
    .IA(\IDLY/$1I328/M01 ),
    .IB(\IDLY/$1I328/M23 ),
    .O(IRDY_M),
    .SEL(CFG246)
  );
  X_OR2   \IDLY/$1I328/M01/$1I38  (
    .I0(\IDLY/$1I328/M01/M1 ),
    .I1(\IDLY/$1I328/M01/M0 ),
    .O(\IDLY/$1I328/M01 )
  );
  X_AND3   \IDLY/$1I328/M01/$1I31  (
    .I0(\NlwInverterSignal_IDLY/$1I328/M01/$1I31/I0 ),
    .I1(\IDLY/$1N332 ),
    .I2(IRDY_I),
    .O(\IDLY/$1I328/M01/M0 )
  );
  X_AND3   \IDLY/$1I328/M01/$1I30  (
    .I0(\IDLY/D3_4180 ),
    .I1(\IDLY/$1N332 ),
    .I2(CFG245),
    .O(\IDLY/$1I328/M01/M1 )
  );
  X_OR2   \IDLY/$1I328/M23/$1I38  (
    .I0(\IDLY/$1I328/M23/M1 ),
    .I1(\IDLY/$1I328/M23/M0 ),
    .O(\IDLY/$1I328/M23 )
  );
  X_AND3   \IDLY/$1I328/M23/$1I31  (
    .I0(\NlwInverterSignal_IDLY/$1I328/M23/$1I31/I0 ),
    .I1(\IDLY/$1N332 ),
    .I2(\IDLY/D4_4181 ),
    .O(\IDLY/$1I328/M23/M0 )
  );
  X_AND3   \IDLY/$1I328/M23/$1I30  (
    .I0(\IDLY/D5_4182 ),
    .I1(\IDLY/$1N332 ),
    .I2(CFG245),
    .O(\IDLY/$1I328/M23/M1 )
  );
  X_ONE   \IDLY/$1I331/$1I2220  (
    .O(\IDLY/$1I331/$1N2216 )
  );
  X_BUF   \IDLY/$1I331/H  (
    .I(\IDLY/$1I331/$1N2216 ),
    .O(\IDLY/$1N332 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \DATA_VLD/SDV_FF  (
    .CE(VCC),
    .CLK(CLK),
    .I(\DATA_VLD/NS_SDV ),
    .O(S_DATA_VLD),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND3   \DATA_VLD/$1I426  (
    .I0(\NlwInverterSignal_DATA_VLD/$1I426/I0 ),
    .I1(\NlwInverterSignal_DATA_VLD/$1I426/I1 ),
    .I2(S_DATA_INT),
    .O(\DATA_VLD/NS_SDV )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \DATA_VLD/MDV_FF  (
    .CE(VCC),
    .CLK(CLK),
    .I(\DATA_VLD/NS_MDV ),
    .O(M_DATA_VLD),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND3   \DATA_VLD/$1I328  (
    .I0(\NlwInverterSignal_DATA_VLD/$1I328/I0 ),
    .I1(\NlwInverterSignal_DATA_VLD/$1I328/I1 ),
    .I2(M_DATA_INT),
    .O(\DATA_VLD/NS_MDV )
  );
  X_AND3   \SRC_EN/$1I742  (
    .I0(\NlwInverterSignal_SRC_EN/$1I742/I0 ),
    .I1(M_WRDN),
    .I2(\SRC_EN/MDATA_EQN ),
    .O(NlwRenamedSig_OI_M_SRC_EN)
  );
  X_AND2   \SRC_EN/$1I656  (
    .I0(\NlwInverterSignal_SRC_EN/$1I656/I0 ),
    .I1(\SRC_EN/S_SRC_PRE ),
    .O(S_SRC_EN)
  );
  X_AND4   \SRC_EN/$1I615  (
    .I0(\NlwInverterSignal_SRC_EN/$1I615/I0 ),
    .I1(NEWDATA),
    .I2(M_READY),
    .I3(M_DATA_INT),
    .O(\SRC_EN/MDATA_EQN )
  );
  X_AND3   \SRC_EN/$1I570  (
    .I0(S_DATA_INT),
    .I1(S_FIRST),
    .I2(S_READY),
    .O(\SRC_EN/SFIRST_EQN )
  );
  X_OR2   \SRC_EN/$1I565  (
    .I0(\SRC_EN/SDATA_EQN ),
    .I1(\SRC_EN/SFIRST_EQN ),
    .O(\SRC_EN/S_SRC_PRE )
  );
  X_AND4   \SRC_EN/$1I558  (
    .I0(\NlwInverterSignal_SRC_EN/$1I558/I0 ),
    .I1(\TSTOP_I- ),
    .I2(NEWDATA),
    .I3(S_READY),
    .O(\SRC_EN/SDATA_EQN )
  );
  X_BUF   \SRC_EN/$1I736/NC  (
    .I(CLK),
    .O(\NLW_SRC_EN/$1I736/NC_O_UNCONNECTED )
  );
  X_BUF   \SRC_EN/$1I737/NC  (
    .I(NlwRenamedSig_OI_RST),
    .O(\NLW_SRC_EN/$1I737/NC_O_UNCONNECTED )
  );
  X_OR2   \OUT_CE/$3I1093  (
    .I0(\OUT_CE/$3N1090 ),
    .I1(\OUT_CE/$3N1089 ),
    .O(\OUT_CE/FIRST )
  );
  X_AND2   \OUT_CE/$3I1092  (
    .I0(S_FIRST),
    .I1(S_DATA_INT),
    .O(\OUT_CE/$3N1089 )
  );
  X_AND2   \OUT_CE/$3I1091  (
    .I0(M_FIRST),
    .I1(M_DATA_INT),
    .O(\OUT_CE/$3N1090 )
  );
  X_AND2   \OUT_CE/$3I1079  (
    .I0(\NlwInverterSignal_OUT_CE/$3I1079/I0 ),
    .I1(M_DATA_INT),
    .O(\NlwInverterSignal_OUT_CE/$3I1079/O )
  );
  X_AND2   \OUT_CE/$3I1078  (
    .I0(\NlwInverterSignal_OUT_CE/$3I1078/I0 ),
    .I1(S_DATA_INT),
    .O(\NlwInverterSignal_OUT_CE/$3I1078/O )
  );
  X_OR3   \OUT_CE/$3I1067  (
    .I0(ADDR_BE),
    .I1(\OUT_CE/FIRST ),
    .I2(FAIL64_INT),
    .O(\OUT_CE/FFA_4285 )
  );
  X_AND3   \OUT_CE/$3I1062  (
    .I0(\NlwInverterSignal_OUT_CE/$3I1062/I0 ),
    .I1(\NlwInverterSignal_OUT_CE/$3I1062/I1 ),
    .I2(M_DATA_INT),
    .O(\OUT_CE/MND_4275 )
  );
  X_AND3   \OUT_CE/$3I1061  (
    .I0(\NlwInverterSignal_OUT_CE/$3I1061/I0 ),
    .I1(\NlwInverterSignal_OUT_CE/$3I1061/I1 ),
    .I2(S_DATA_INT),
    .O(\OUT_CE/SND_4267 )
  );
  X_OR2   \OUT_CE/$3I1057  (
    .I0(ADDR_BE),
    .I1(\OUT_CE/FIRST ),
    .O(\OUT_CE/$3N1041 )
  );
  X_AND2   \OUT_CE/$3I1056  (
    .I0(\NlwInverterSignal_OUT_CE/$3I1056/I0 ),
    .I1(\OUT_CE/$3N1041 ),
    .O(\OUT_CE/FANF_4266 )
  );
  X_AND2   \OUT_CE/$2I1086  (
    .I0(\NlwInverterSignal_OUT_CE/$2I1086/I0 ),
    .I1(\NlwInverterSignal_OUT_CE/$2I1086/I1 ),
    .O(\OUT_CE/M_CE_XX1 )
  );
  X_AND2   \OUT_CE/$2I1085  (
    .I0(\NlwInverterSignal_OUT_CE/$2I1085/I0 ),
    .I1(\NlwInverterSignal_OUT_CE/$2I1085/I1 ),
    .O(\OUT_CE/M_CE_XX0 )
  );
  X_AND2   \OUT_CE/$2I1084  (
    .I0(\NlwInverterSignal_OUT_CE/$2I1084/I0 ),
    .I1(\NlwInverterSignal_OUT_CE/$2I1084/I1 ),
    .O(\OUT_CE/S_CE_XX1 )
  );
  X_AND2   \OUT_CE/$2I1083  (
    .I0(\NlwInverterSignal_OUT_CE/$2I1083/I0 ),
    .I1(\NlwInverterSignal_OUT_CE/$2I1083/I1 ),
    .O(\OUT_CE/S_CE_XX0 )
  );
  X_MUX2   \OUT_CE/$2I1053  (
    .IA(\OUT_CE/SOFT_CE0 ),
    .IB(\OUT_CE/SOFT_CE1 ),
    .O(\OUT_CE/SOFT_CE ),
    .SEL(IRDY_F)
  );
  X_OR3   \OUT_CE/$2I1052  (
    .I0(\OUT_CE/S_CE_XX0 ),
    .I1(\OUT_CE/FFA_4285 ),
    .I2(\OUT_CE/M_CE_XX0 ),
    .O(\OUT_CE/SOFT_CE0 )
  );
  X_OR3   \OUT_CE/$2I1051  (
    .I0(\OUT_CE/S_CE_XX1 ),
    .I1(\OUT_CE/FFA_4285 ),
    .I2(\OUT_CE/M_CE_XX1 ),
    .O(\OUT_CE/SOFT_CE1 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \OUT_CE/PAR_CE  (
    .CE(VCC),
    .CLK(CLK),
    .I(\OUT_CE/NS_PAR_CE ),
    .O(PAR_CE),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_OR3   \OUT_CE/$2I1016  (
    .I0(\OUT_CE/S_CE_P1 ),
    .I1(\OUT_CE/FFA_4285 ),
    .I2(\OUT_CE/M_CE_P1 ),
    .O(\OUT_CE/NS_PAR_CE1 )
  );
  X_AND2   \OUT_CE/$2I1015  (
    .I0(\NlwInverterSignal_OUT_CE/$2I1015/I0 ),
    .I1(\NlwInverterSignal_OUT_CE/$2I1015/I1 ),
    .O(\OUT_CE/M_CE_P1 )
  );
  X_AND2   \OUT_CE/$2I1013  (
    .I0(\NlwInverterSignal_OUT_CE/$2I1013/I0 ),
    .I1(\NlwInverterSignal_OUT_CE/$2I1013/I1 ),
    .O(\OUT_CE/M_CE_P0 )
  );
  X_AND2   \OUT_CE/$2I1012  (
    .I0(\NlwInverterSignal_OUT_CE/$2I1012/I0 ),
    .I1(\NlwInverterSignal_OUT_CE/$2I1012/I1 ),
    .O(\OUT_CE/S_CE_P0 )
  );
  X_OR3   \OUT_CE/$2I1011  (
    .I0(\OUT_CE/S_CE_P0 ),
    .I1(\OUT_CE/FFA_4285 ),
    .I2(\OUT_CE/M_CE_P0 ),
    .O(\OUT_CE/NS_PAR_CE0 )
  );
  X_MUX2   \OUT_CE/$2I1008  (
    .IA(\OUT_CE/NS_PAR_CE0 ),
    .IB(\OUT_CE/NS_PAR_CE1 ),
    .O(\OUT_CE/NS_PAR_CE ),
    .SEL(IRDY_M)
  );
  X_AND2   \OUT_CE/$2I1007  (
    .I0(\NlwInverterSignal_OUT_CE/$2I1007/I0 ),
    .I1(\NlwInverterSignal_OUT_CE/$2I1007/I1 ),
    .O(\OUT_CE/S_CE_P1 )
  );
  X_AND2   \OUT_CE/$1I980  (
    .I0(\NlwInverterSignal_OUT_CE/$1I980/I0 ),
    .I1(\OUT_CE/SND_4267 ),
    .O(\OUT_CE/S_ND_T1 )
  );
  X_MUX2   \OUT_CE/$1I979  (
    .IA(\OUT_CE/ZERO_ND_T0 ),
    .IB(\OUT_CE/ZERO_ND_T1 ),
    .O(\OUT_CE/NS_NEWDATA ),
    .SEL(TRDY_M)
  );
  X_OR3   \OUT_CE/$1I977  (
    .I0(\OUT_CE/S_ND_T0 ),
    .I1(\OUT_CE/FANF_4266 ),
    .I2(\OUT_CE/M_ND_T0 ),
    .O(\OUT_CE/ZERO_ND_T0 )
  );
  X_AND2   \OUT_CE/$1I976  (
    .I0(\NlwInverterSignal_OUT_CE/$1I976/I0 ),
    .I1(\OUT_CE/SND_4267 ),
    .O(\OUT_CE/S_ND_T0 )
  );
  X_AND2   \OUT_CE/$1I975  (
    .I0(\NlwInverterSignal_OUT_CE/$1I975/I0 ),
    .I1(\OUT_CE/MND_4275 ),
    .O(\OUT_CE/M_ND_T0 )
  );
  X_AND2   \OUT_CE/$1I972  (
    .I0(\NlwInverterSignal_OUT_CE/$1I972/I0 ),
    .I1(\OUT_CE/MND_4275 ),
    .O(\OUT_CE/M_ND_T1 )
  );
  X_OR3   \OUT_CE/$1I971  (
    .I0(\OUT_CE/S_ND_T1 ),
    .I1(\OUT_CE/FANF_4266 ),
    .I2(\OUT_CE/M_ND_T1 ),
    .O(\OUT_CE/ZERO_ND_T1 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \OUT_CE/NDFF  (
    .CE(VCC),
    .CLK(CLK),
    .I(\OUT_CE/NS_NEWDATA ),
    .O(NEWDATA),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_ZERO   \OUT_CE/$1I987/$1I2218  (
    .O(\OUT_CE/$1I987/$1N2216 )
  );
  X_BUF   \OUT_CE/$1I987/L  (
    .I(\OUT_CE/$1I987/$1N2216 ),
    .O(\OUT_CE/$1N989 )
  );
  X_ONE   \OUT_CE/$1I988/$1I2220  (
    .O(\OUT_CE/$1I988/$1N2216 )
  );
  X_BUF   \OUT_CE/$1I988/H  (
    .I(\OUT_CE/$1I988/$1N2216 ),
    .O(\OUT_CE/$1N968 )
  );
  X_ZERO   \OUT_CE/$2I1022/$1I2218  (
    .O(\OUT_CE/$2I1022/$1N2216 )
  );
  X_BUF   \OUT_CE/$2I1022/L  (
    .I(\OUT_CE/$2I1022/$1N2216 ),
    .O(\OUT_CE/$2N1025 )
  );
  X_ONE   \OUT_CE/$2I1023/$1I2220  (
    .O(\OUT_CE/$2I1023/$1N2216 )
  );
  X_BUF   \OUT_CE/$2I1023/H  (
    .I(\OUT_CE/$2I1023/$1N2216 ),
    .O(\OUT_CE/$2N1024 )
  );
  X_ONE   \OUT_CE/$2I1049/$1I2220  (
    .O(\OUT_CE/$2I1049/$1N2216 )
  );
  X_BUF   \OUT_CE/$2I1049/H  (
    .I(\OUT_CE/$2I1049/$1N2216 ),
    .O(\OUT_CE/$2N1067 )
  );
  X_ZERO   \OUT_CE/$2I1050/$1I2218  (
    .O(\OUT_CE/$2I1050/$1N2216 )
  );
  X_BUF   \OUT_CE/$2I1050/L  (
    .I(\OUT_CE/$2I1050/$1N2216 ),
    .O(\OUT_CE/$2N1066 )
  );
  X_AND3   \OUT_CE/MAGICBOX/PCI_CE  (
    .I0(\NlwInverterSignal_OUT_CE/MAGICBOX/PCI_CE/I0 ),
    .I1(\OUT_CE/MAGICBOX/I1_NAND_IRDY_4238 ),
    .I2(\OUT_CE/MAGICBOX/I3_NAND_TRDY_4239 ),
    .O(\NlwInverterSignal_OUT_CE/MAGICBOX/PCI_CE/O )
  );
  X_AND2   \OUT_CE/MAGICBOX/I3_NAND_TRDY  (
    .I0(\NlwInverterSignal_OUT_CE/MAGICBOX/I3_NAND_TRDY/I0 ),
    .I1(\NlwInverterSignal_OUT_CE/MAGICBOX/I3_NAND_TRDY/I1 ),
    .O(\NlwInverterSignal_OUT_CE/MAGICBOX/I3_NAND_TRDY/O )
  );
  X_AND2   \OUT_CE/MAGICBOX/I1_NAND_IRDY  (
    .I0(\NlwInverterSignal_OUT_CE/MAGICBOX/I1_NAND_IRDY/I0 ),
    .I1(\NlwInverterSignal_OUT_CE/MAGICBOX/I1_NAND_IRDY/I1 ),
    .O(\NlwInverterSignal_OUT_CE/MAGICBOX/I1_NAND_IRDY/O )
  );
  X_AND2   \OUT_CE/$4I1005/$1I9  (
    .I0(\OUT_CE/SOFT_CE ),
    .I1(CFG251),
    .O(\OUT_CE/$4I1005/M1 )
  );
  X_OR2   \OUT_CE/$4I1005/$1I8  (
    .I0(\OUT_CE/$4I1005/M1 ),
    .I1(\OUT_CE/$4I1005/M0 ),
    .O(PCI_CE)
  );
  X_AND2   \OUT_CE/$4I1005/$1I7  (
    .I0(\NlwInverterSignal_OUT_CE/$4I1005/$1I7/I0 ),
    .I1(\OUT_CE/HARD_CE ),
    .O(\OUT_CE/$4I1005/M0 )
  );
  X_AND2   \OUT_SEL/$1I952  (
    .I0(\OUT_SEL/S_IN ),
    .I1(IRDY_M),
    .O(\OUT_SEL/$1N959 )
  );
  X_OR2   \OUT_SEL/$1I951  (
    .I0(\OUT_SEL/$1N959 ),
    .I1(\OUT_SEL/$1N958 ),
    .O(\OUT_SEL/SEL64_IN )
  );
  X_AND2   \OUT_SEL/$1I940  (
    .I0(TRDY_M),
    .I1(\OUT_SEL/M_IN ),
    .O(\OUT_SEL/$1N958 )
  );
  X_AND3   \OUT_SEL/$1I916  (
    .I0(\NlwInverterSignal_OUT_SEL/$1I916/I0 ),
    .I1(\NlwInverterSignal_OUT_SEL/$1I916/I1 ),
    .I2(S_DATA_INT),
    .O(\OUT_SEL/S_IN )
  );
  X_AND4   \OUT_SEL/$1I913  (
    .I0(\NlwInverterSignal_OUT_SEL/$1I913/I0 ),
    .I1(\NlwInverterSignal_OUT_SEL/$1I913/I1 ),
    .I2(\NlwInverterSignal_OUT_SEL/$1I913/I2 ),
    .I3(M_DATA_INT),
    .O(\OUT_SEL/M_IN )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \OUT_SEL/OSEL64_FF  (
    .CE(VCC),
    .CLK(CLK),
    .I(\OUT_SEL/SEL64_IN ),
    .O(OUT_SEL64),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND2   \OUT_SEL/$1I897  (
    .I0(\NlwInverterSignal_OUT_SEL/$1I897/I0 ),
    .I1(S_DATA_INT),
    .O(\OUT_SEL/$1N898 )
  );
  X_OR2   \OUT_SEL/$1I896  (
    .I0(M_DATA_INT),
    .I1(\OUT_SEL/$1N898 ),
    .O(\OUT_SEL/$1N851 )
  );
  X_AND2   \OUT_SEL/$1I853  (
    .I0(\NlwInverterSignal_OUT_SEL/$1I853/I0 ),
    .I1(\OUT_SEL/$1N765 ),
    .O(SHADOW_CE64)
  );
  X_AND2   \OUT_SEL/$1I849  (
    .I0(\NlwInverterSignal_OUT_SEL/$1I849/I0 ),
    .I1(\OUT_SEL/$1N851 ),
    .O(SHADOW_CE)
  );
  X_AND2   \OUT_SEL/$1I836  (
    .I0(\OUT_SEL/S_IN ),
    .I1(IRDY_M),
    .O(\OUT_SEL/$1N821 )
  );
  X_AND2   \OUT_SEL/$1I815  (
    .I0(TRDY_M),
    .I1(\OUT_SEL/M_IN ),
    .O(\OUT_SEL/$1N826 )
  );
  X_OR2   \OUT_SEL/$1I814  (
    .I0(\OUT_SEL/$1N821 ),
    .I1(\OUT_SEL/$1N826 ),
    .O(\OUT_SEL/SEL_IN )
  );
  X_OR2   \OUT_SEL/$1I767  (
    .I0(M_DATA_INT),
    .I1(\OUT_SEL/$1N766 ),
    .O(\OUT_SEL/$1N765 )
  );
  X_AND2   \OUT_SEL/$1I758  (
    .I0(\NlwInverterSignal_OUT_SEL/$1I758/I0 ),
    .I1(S_DATA_INT),
    .O(\OUT_SEL/$1N766 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \OUT_SEL/OSEL_FF  (
    .CE(VCC),
    .CLK(CLK),
    .I(\OUT_SEL/SEL_IN ),
    .O(OUT_SEL),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND4   \ADDR_VLD/$1I4008  (
    .I0(\NlwInverterSignal_ADDR_VLD/$1I4008/I0 ),
    .I1(\NlwInverterSignal_ADDR_VLD/$1I4008/I1 ),
    .I2(\ADDR_VLD/TEMP_1 ),
    .I3(\ADDR_VLD/TEMP_2 ),
    .O(ADDR_VLD64)
  );
  X_AND2   \ADDR_VLD/$1I4005  (
    .I0(\NlwInverterSignal_ADDR_VLD/$1I4005/I0 ),
    .I1(M_DATA_INT),
    .O(\NlwInverterSignal_ADDR_VLD/$1I4005/O )
  );
  X_AND3   \ADDR_VLD/$1I4000  (
    .I0(SLOT64),
    .I1(\ADDR_VLD/REQ64Q- ),
    .I2(\ADDR_VLD/FRAMEQ- ),
    .O(\ADDR_VLD/TEMP_1 )
  );
  X_AND2   \ADDR_VLD/$1I3989  (
    .I0(\NlwInverterSignal_ADDR_VLD/$1I3989/I0 ),
    .I1(M_DATA_INT),
    .O(\NlwInverterSignal_ADDR_VLD/$1I3989/O )
  );
  X_AND2   \ADDR_VLD/$1I3986  (
    .I0(\NlwInverterSignal_ADDR_VLD/$1I3986/I0 ),
    .I1(M_DATA_INT),
    .O(\NlwInverterSignal_ADDR_VLD/$1I3986/O )
  );
  X_AND2   \ADDR_VLD/$1I3983  (
    .I0(\NlwInverterSignal_ADDR_VLD/$1I3983/I0 ),
    .I1(M_DATA_INT),
    .O(\NlwInverterSignal_ADDR_VLD/$1I3983/O )
  );
  X_AND2   \ADDR_VLD/$1I3980  (
    .I0(\NlwInverterSignal_ADDR_VLD/$1I3980/I0 ),
    .I1(M_DATA_INT),
    .O(\NlwInverterSignal_ADDR_VLD/$1I3980/O )
  );
  X_AND2   \ADDR_VLD/$1I3967  (
    .I0(\ADDR_VLD/FRAMEQ- ),
    .I1(IDSEL),
    .O(\ADDR_VLD/TEMP_0 )
  );
  X_AND3   \ADDR_VLD/$1I3963  (
    .I0(\NlwInverterSignal_ADDR_VLD/$1I3963/I0 ),
    .I1(\ADDR_VLD/TEMP_0 ),
    .I2(\ADDR_VLD/$1N3964 ),
    .O(NlwRenamedSig_OI_CFG_VLD)
  );
  X_AND3   \ADDR_VLD/$1I3894  (
    .I0(\NlwInverterSignal_ADDR_VLD/$1I3894/I0 ),
    .I1(\ADDR_VLD/FRAMEQ- ),
    .I2(\ADDR_VLD/$1N3898 ),
    .O(ADDR_VLD1)
  );
  X_AND3   \ADDR_VLD/$1I3880  (
    .I0(\NlwInverterSignal_ADDR_VLD/$1I3880/I0 ),
    .I1(\ADDR_VLD/FRAMEQ- ),
    .I2(\ADDR_VLD/$1N3884 ),
    .O(ADDR_VLD0)
  );
  X_AND3   \ADDR_VLD/$1I3867  (
    .I0(\NlwInverterSignal_ADDR_VLD/$1I3867/I0 ),
    .I1(\ADDR_VLD/FRAMEQ- ),
    .I2(\ADDR_VLD/$1N3858 ),
    .O(NlwRenamedSig_OI_ADDR_VLD)
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \ADDR_VLD/$1I3821  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(CLK),
    .I(\FRAME- ),
    .O(\ADDR_VLD/FRAMEQ- ),
    .RST(GND)
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \ADDR_VLD/$1I3811  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(CLK),
    .I(\REQ64- ),
    .O(\ADDR_VLD/REQ64Q- ),
    .RST(GND)
  );
  X_AND2   \EOT/$1I619  (
    .I0(\EOT/$1N631 ),
    .I1(\EOT/EQN-V1 ),
    .O(\EOT/$1N630 )
  );
  X_OR2   \EOT/$1I618  (
    .I0(\EOT/$1N630 ),
    .I1(\EOT/EQN-W1 ),
    .O(\EOT/NS_1 )
  );
  X_OR2   \EOT/$1I617  (
    .I0(\NlwInverterSignal_EOT/$1I617/I0 ),
    .I1(\NlwInverterSignal_EOT/$1I617/I1 ),
    .O(\EOT/$1N631 )
  );
  X_AND2   \EOT/$1I616  (
    .I0(\NlwInverterSignal_EOT/$1I616/I0 ),
    .I1(EOT),
    .O(\EOT/$1N627 )
  );
  X_OR2   \EOT/$1I615  (
    .I0(\NlwInverterSignal_EOT/$1I615/I0 ),
    .I1(\NlwInverterSignal_EOT/$1I615/I1 ),
    .O(\EOT/$1N624 )
  );
  X_AND2   \EOT/$1I614  (
    .I0(\IFRAME_I- ),
    .I1(M_DATA_INT),
    .O(\EOT/EQN-V1 )
  );
  X_OR2   \EOT/$1I613  (
    .I0(\EOT/$1N623 ),
    .I1(\EOT/$1N627 ),
    .O(\EOT/EQN-W1 )
  );
  X_AND2   \EOT/$1I610  (
    .I0(\EOT/$1N624 ),
    .I1(S_DATA_INT),
    .O(\EOT/$1N623 )
  );
  X_AND2   \EOT/$1I591  (
    .I0(\EOT/$1N603 ),
    .I1(\EOT/EQN-V0 ),
    .O(\EOT/$1N658 )
  );
  X_OR2   \EOT/$1I590  (
    .I0(\EOT/$1N658 ),
    .I1(\EOT/EQN-W0 ),
    .O(\EOT/NS_0 )
  );
  X_OR2   \EOT/$1I589  (
    .I0(\NlwInverterSignal_EOT/$1I589/I0 ),
    .I1(\NlwInverterSignal_EOT/$1I589/I1 ),
    .O(\EOT/$1N603 )
  );
  X_AND2   \EOT/$1I588  (
    .I0(\NlwInverterSignal_EOT/$1I588/I0 ),
    .I1(EOT),
    .O(\EOT/EQN-W0 )
  );
  X_AND2   \EOT/$1I585  (
    .I0(\IFRAME_I- ),
    .I1(M_DATA_INT),
    .O(\EOT/EQN-V0 )
  );
  X_MUX2   \EOT/$1I579  (
    .IA(\EOT/NS_0 ),
    .IB(\EOT/NS_1 ),
    .O(\EOT/EOT_D ),
    .SEL(FRAME_I)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \EOT/EOT_DL  (
    .CE(VCC),
    .CLK(CLK),
    .I(EOT),
    .O(\EOT/EOT_DL_4369 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \EOT/EOT_FF  (
    .CE(VCC),
    .CLK(CLK),
    .I(\EOT/EOT_D ),
    .O(EOT),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR4   \PCI-PAR/$7I3007  (
    .I0(CBE_I0),
    .I1(CBE_I1),
    .I2(CBE_I2),
    .I3(CBE_I3),
    .O(\PCI-PAR/PREP )
  );
  X_MUX2   \PCI-PAR/$7I3006  (
    .IA(\PCI-PAR/PREP ),
    .IB(\PCI-PAR/PREN ),
    .O(NS_PAR),
    .SEL(\PCI-PAR/AD_PAR )
  );
  X_XOR4   \PCI-PAR/$7I2985  (
    .I0(CBE_I0),
    .I1(CBE_I1),
    .I2(CBE_I2),
    .I3(CBE_I3),
    .O(\NlwInverterSignal_PCI-PAR/$7I2985/O )
  );
  X_XOR4   \PCI-PAR/$7I2974  (
    .I0(CBE_I4),
    .I1(CBE_I5),
    .I2(CBE_I6),
    .I3(CBE_I7),
    .O(\NlwInverterSignal_PCI-PAR/$7I2974/O )
  );
  X_MUX2   \PCI-PAR/$7I2973  (
    .IA(\PCI-PAR/PRE64P ),
    .IB(\PCI-PAR/PRE64N ),
    .O(NS_PAR64),
    .SEL(\PCI-PAR/AD_PAR64 )
  );
  X_XOR4   \PCI-PAR/$7I2972  (
    .I0(CBE_I4),
    .I1(CBE_I5),
    .I2(CBE_I6),
    .I3(CBE_I7),
    .O(\PCI-PAR/PRE64P )
  );
  X_XOR2   \PCI-PAR/X46  (
    .I0(\PCI-PAR/X14O ),
    .I1(\PCI-PAR/X15O ),
    .O(\PCI-PAR/P7O )
  );
  X_XOR2   \PCI-PAR/X43  (
    .I0(\PCI-PAR/X12O ),
    .I1(\PCI-PAR/X13O ),
    .O(\PCI-PAR/P6O )
  );
  X_XOR2   \PCI-PAR/X40  (
    .I0(\PCI-PAR/X10O ),
    .I1(\PCI-PAR/X11O ),
    .O(\PCI-PAR/P5O )
  );
  X_XOR2   \PCI-PAR/X37  (
    .I0(\PCI-PAR/X8O ),
    .I1(\PCI-PAR/X9O ),
    .O(\PCI-PAR/P4O )
  );
  X_XOR4   \PCI-PAR/X45  (
    .I0(\PCI-PAR/DOQ56 ),
    .I1(\PCI-PAR/DOQ57 ),
    .I2(\PCI-PAR/DOQ58 ),
    .I3(\PCI-PAR/DOQ59 ),
    .O(\PCI-PAR/X14O )
  );
  X_XOR4   \PCI-PAR/X44  (
    .I0(\PCI-PAR/DOQ52 ),
    .I1(\PCI-PAR/DOQ53 ),
    .I2(\PCI-PAR/DOQ54 ),
    .I3(\PCI-PAR/DOQ55 ),
    .O(\PCI-PAR/X13O )
  );
  X_XOR4   \PCI-PAR/X42  (
    .I0(\PCI-PAR/DOQ48 ),
    .I1(\PCI-PAR/DOQ49 ),
    .I2(\PCI-PAR/DOQ50 ),
    .I3(\PCI-PAR/DOQ51 ),
    .O(\PCI-PAR/X12O )
  );
  X_XOR4   \PCI-PAR/X41  (
    .I0(\PCI-PAR/DOQ44 ),
    .I1(\PCI-PAR/DOQ45 ),
    .I2(\PCI-PAR/DOQ46 ),
    .I3(\PCI-PAR/DOQ47 ),
    .O(\PCI-PAR/X11O )
  );
  X_XOR4   \PCI-PAR/X39  (
    .I0(\PCI-PAR/DOQ40 ),
    .I1(\PCI-PAR/DOQ41 ),
    .I2(\PCI-PAR/DOQ42 ),
    .I3(\PCI-PAR/DOQ43 ),
    .O(\PCI-PAR/X10O )
  );
  X_XOR4   \PCI-PAR/X38  (
    .I0(\PCI-PAR/DOQ36 ),
    .I1(\PCI-PAR/DOQ37 ),
    .I2(\PCI-PAR/DOQ38 ),
    .I3(\PCI-PAR/DOQ39 ),
    .O(\PCI-PAR/X9O )
  );
  X_XOR4   \PCI-PAR/X36  (
    .I0(\PCI-PAR/DOQ32 ),
    .I1(\PCI-PAR/DOQ33 ),
    .I2(\PCI-PAR/DOQ34 ),
    .I3(\PCI-PAR/DOQ35 ),
    .O(\PCI-PAR/X8O )
  );
  X_XOR4   \PCI-PAR/X47  (
    .I0(\PCI-PAR/DOQ60 ),
    .I1(\PCI-PAR/DOQ61 ),
    .I2(\PCI-PAR/DOQ62 ),
    .I3(\PCI-PAR/DOQ63 ),
    .O(\PCI-PAR/X15O )
  );
  X_XOR4   \PCI-PAR/$6I3192  (
    .I0(\PCI-PAR/P4O ),
    .I1(\PCI-PAR/P5O ),
    .I2(\PCI-PAR/P6O ),
    .I3(\PCI-PAR/P7O ),
    .O(\PCI-PAR/AD_PAR64 )
  );
  X_XOR2   \PCI-PAR/X25  (
    .I0(\PCI-PAR/X0O ),
    .I1(\PCI-PAR/X1O ),
    .O(\PCI-PAR/P0O )
  );
  X_XOR2   \PCI-PAR/X28  (
    .I0(\PCI-PAR/X2O ),
    .I1(\PCI-PAR/X3O ),
    .O(\PCI-PAR/P1O )
  );
  X_XOR2   \PCI-PAR/X31  (
    .I0(\PCI-PAR/X4O ),
    .I1(\PCI-PAR/X5O ),
    .O(\PCI-PAR/P2O )
  );
  X_XOR2   \PCI-PAR/X34  (
    .I0(\PCI-PAR/X6O ),
    .I1(\PCI-PAR/X7O ),
    .O(\PCI-PAR/P3O )
  );
  X_XOR4   \PCI-PAR/$5I3093  (
    .I0(\PCI-PAR/P0O ),
    .I1(\PCI-PAR/P1O ),
    .I2(\PCI-PAR/P2O ),
    .I3(\PCI-PAR/P3O ),
    .O(\PCI-PAR/AD_PAR )
  );
  X_XOR4   \PCI-PAR/X35  (
    .I0(\PCI-PAR/DOQ28 ),
    .I1(\PCI-PAR/DOQ29 ),
    .I2(\PCI-PAR/DOQ30 ),
    .I3(\PCI-PAR/DOQ31 ),
    .O(\PCI-PAR/X7O )
  );
  X_XOR4   \PCI-PAR/X33  (
    .I0(\PCI-PAR/DOQ24 ),
    .I1(\PCI-PAR/DOQ25 ),
    .I2(\PCI-PAR/DOQ26 ),
    .I3(\PCI-PAR/DOQ27 ),
    .O(\PCI-PAR/X6O )
  );
  X_XOR4   \PCI-PAR/X32  (
    .I0(\PCI-PAR/DOQ20 ),
    .I1(\PCI-PAR/DOQ21 ),
    .I2(\PCI-PAR/DOQ22 ),
    .I3(\PCI-PAR/DOQ23 ),
    .O(\PCI-PAR/X5O )
  );
  X_XOR4   \PCI-PAR/X30  (
    .I0(\PCI-PAR/DOQ16 ),
    .I1(\PCI-PAR/DOQ17 ),
    .I2(\PCI-PAR/DOQ18 ),
    .I3(\PCI-PAR/DOQ19 ),
    .O(\PCI-PAR/X4O )
  );
  X_XOR4   \PCI-PAR/X29  (
    .I0(\PCI-PAR/DOQ12 ),
    .I1(\PCI-PAR/DOQ13 ),
    .I2(\PCI-PAR/DOQ14 ),
    .I3(\PCI-PAR/DOQ15 ),
    .O(\PCI-PAR/X3O )
  );
  X_XOR4   \PCI-PAR/X27  (
    .I0(\PCI-PAR/DOQ8 ),
    .I1(\PCI-PAR/DOQ9 ),
    .I2(\PCI-PAR/DOQ10 ),
    .I3(\PCI-PAR/DOQ11 ),
    .O(\PCI-PAR/X2O )
  );
  X_XOR4   \PCI-PAR/X26  (
    .I0(\PCI-PAR/DOQ4 ),
    .I1(\PCI-PAR/DOQ5 ),
    .I2(\PCI-PAR/DOQ6 ),
    .I3(\PCI-PAR/DOQ7 ),
    .O(\PCI-PAR/X1O )
  );
  X_XOR4   \PCI-PAR/X24  (
    .I0(\PCI-PAR/DOQ0 ),
    .I1(\PCI-PAR/DOQ1 ),
    .I2(\PCI-PAR/DOQ2 ),
    .I3(\PCI-PAR/DOQ3 ),
    .O(\PCI-PAR/X0O )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-PAR/APERR_N  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(CLK),
    .I(\PCI-PAR/PRE_APERR_N ),
    .O(APERR_N),
    .RST(GND)
  );
  X_AND2   \PCI-PAR/$4I3163  (
    .I0(PERR_EN),
    .I1(ADDR_VLD64),
    .O(\PCI-PAR/CHECK64 )
  );
  X_AND2   \PCI-PAR/$4I3157  (
    .I0(PERR_EN),
    .I1(ADDR_VLD1),
    .O(\PCI-PAR/CHECK32 )
  );
  X_MUX2   \PCI-PAR/$4I3133  (
    .IA(\PCI-PAR/PAP_0 ),
    .IB(\PCI-PAR/PAP_1 ),
    .O(\PCI-PAR/PRE_APERR_N ),
    .SEL(PAR64_I)
  );
  X_XOR2   \PCI-PAR/$4I3131  (
    .I0(\PCI-PAR/PER64_4858 ),
    .I1(\PCI-PAR/$4N3107 ),
    .O(\PCI-PAR/$4N3110 )
  );
  X_XOR2   \PCI-PAR/$4I3128  (
    .I0(\PCI-PAR/PER64_4858 ),
    .I1(\PCI-PAR/$4N3125 ),
    .O(\PCI-PAR/$4N3113 )
  );
  X_OR2   \PCI-PAR/$4I3127  (
    .I0(\PCI-PAR/PAP64_0 ),
    .I1(\PCI-PAR/PAP32_0 ),
    .O(\NlwInverterSignal_PCI-PAR/$4I3127/O )
  );
  X_AND2   \PCI-PAR/$4I3120  (
    .I0(\PCI-PAR/$4N3098 ),
    .I1(\PCI-PAR/CHECK32 ),
    .O(\PCI-PAR/PAP32_0 )
  );
  X_AND2   \PCI-PAR/$4I3112  (
    .I0(\PCI-PAR/$4N3113 ),
    .I1(\PCI-PAR/CHECK64 ),
    .O(\PCI-PAR/PAP64_0 )
  );
  X_AND2   \PCI-PAR/$4I3111  (
    .I0(\PCI-PAR/$4N3110 ),
    .I1(\PCI-PAR/CHECK64 ),
    .O(\PCI-PAR/PAP64_1 )
  );
  X_AND2   \PCI-PAR/$4I3108  (
    .I0(\PCI-PAR/$4N3109 ),
    .I1(\PCI-PAR/CHECK32 ),
    .O(\PCI-PAR/PAP32_1 )
  );
  X_OR2   \PCI-PAR/$4I3104  (
    .I0(\PCI-PAR/PAP64_1 ),
    .I1(\PCI-PAR/PAP32_1 ),
    .O(\NlwInverterSignal_PCI-PAR/$4I3104/O )
  );
  X_XOR2   \PCI-PAR/$4I3103  (
    .I0(\PCI-PAR/PER_4845 ),
    .I1(PAR_I),
    .O(\PCI-PAR/$4N3109 )
  );
  X_XOR2   \PCI-PAR/$4I3095  (
    .I0(\PCI-PAR/PER_4845 ),
    .I1(PAR_I),
    .O(\PCI-PAR/$4N3098 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$3I3059  (
    .CE(VCC),
    .CLK(CLK),
    .I(M_DATA_INT),
    .O(\PCI-PAR/M_DATAQ ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$3I3058  (
    .CE(VCC),
    .CLK(CLK),
    .I(\PCI-PAR/M_DATAQ ),
    .O(\PCI-PAR/$3N3054 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND3   \PCI-PAR/$3I3057  (
    .I0(\NlwInverterSignal_PCI-PAR/$3I3057/I0 ),
    .I1(PERR_EN),
    .I2(\PCI-PAR/$3N3054 ),
    .O(SET8)
  );
  X_MUX2   \PCI-PAR/$3I3027  (
    .IA(\PCI-PAR/NS_0 ),
    .IB(\PCI-PAR/NS_1 ),
    .O(\NS_PERR- ),
    .SEL(PAR_I)
  );
  X_AND2   \PCI-PAR/$3I3026  (
    .I0(\PCI-PAR/$3N3025 ),
    .I1(\PCI-PAR/PWIN64 ),
    .O(\PCI-PAR/ERR64_1 )
  );
  X_AND2   \PCI-PAR/$3I3023  (
    .I0(\PCI-PAR/$3N3024 ),
    .I1(\PCI-PAR/PWIN ),
    .O(\PCI-PAR/ERR32_1 )
  );
  X_OR2   \PCI-PAR/$3I3018  (
    .I0(\PCI-PAR/ERR64_1 ),
    .I1(\PCI-PAR/ERR32_1 ),
    .O(\NlwInverterSignal_PCI-PAR/$3I3018/O )
  );
  X_XOR2   \PCI-PAR/$3I3017  (
    .I0(\PCI-PAR/PER64_4858 ),
    .I1(PAR64_I),
    .O(\PCI-PAR/$3N3025 )
  );
  X_XOR2   \PCI-PAR/$3I3016  (
    .I0(\PCI-PAR/PER_4845 ),
    .I1(\PCI-PAR/$3N3020 ),
    .O(\PCI-PAR/$3N3024 )
  );
  X_OR3   \PCI-PAR/$3I3005  (
    .I0(IPWIN64),
    .I1(TPWIN64),
    .I2(ADDR_VLD64),
    .O(\PCI-PAR/PWIN64 )
  );
  X_OR3   \PCI-PAR/$3I2999  (
    .I0(IPWIN),
    .I1(TPWIN),
    .I2(ADDR_VLD1),
    .O(\PCI-PAR/PWIN )
  );
  X_OR2   \PCI-PAR/$3I2993  (
    .I0(\PCI-PAR/ERR64_0 ),
    .I1(\PCI-PAR/ERR32_0 ),
    .O(\NlwInverterSignal_PCI-PAR/$3I2993/O )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$3I2944  (
    .CE(VCC),
    .CLK(CLK),
    .I(ADDR_VLD1),
    .O(\PCI-PAR/ADDR_VLDQ ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND2   \PCI-PAR/$3I2940  (
    .I0(PERR_EN),
    .I1(\PCI-PAR/NS_SERR ),
    .O(\NlwInverterSignal_PCI-PAR/$3I2940/O )
  );
  X_INV   \PCI-PAR/$3I2938  (
    .I(\PCI-PAR/NS_OE_SERR ),
    .O(SET14)
  );
  X_OR2   \PCI-PAR/$3I2936  (
    .I0(\NlwInverterSignal_PCI-PAR/$3I2936/I0 ),
    .I1(\PCI-PAR/$3N2935 ),
    .O(\PCI-PAR/NS_OE_SERR )
  );
  X_AND2   \PCI-PAR/$3I2931  (
    .I0(\NlwInverterSignal_PCI-PAR/$3I2931/I0 ),
    .I1(\PCI-PAR/$3N2930 ),
    .O(\PCI-PAR/NS_SERR )
  );
  X_OR2   \PCI-PAR/$3I2929  (
    .I0(NlwRenamedSig_OI_PCI_CMD1),
    .I1(\PCI-PAR/ADDR_VLDQ ),
    .O(\PCI-PAR/$3N2930 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-PAR/OE_SERR_FF  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(CLK),
    .I(\PCI-PAR/NS_OE_SERR ),
    .O(OE_SERR),
    .RST(GND)
  );
  X_AND2   \PCI-PAR/$3I2838  (
    .I0(\PCI-PAR/$3N2766 ),
    .I1(\PCI-PAR/PWIN64 ),
    .O(\PCI-PAR/ERR64_0 )
  );
  X_XOR2   \PCI-PAR/$3I2770  (
    .I0(\PCI-PAR/PER64_4858 ),
    .I1(PAR64_I),
    .O(\PCI-PAR/$3N2766 )
  );
  X_AND2   \PCI-PAR/$3I2764  (
    .I0(\PCI-PAR/$3N2500 ),
    .I1(\PCI-PAR/PWIN ),
    .O(\PCI-PAR/ERR32_0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-PAR/LC_PERR  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .CLK(CLK),
    .I(\NS_PERR- ),
    .O(\PCI-PAR/LC_PERR- ),
    .RST(GND)
  );
  X_INV   \PCI-PAR/$3I2733  (
    .I(\PCI-PAR/LC_PERR- ),
    .O(SET15)
  );
  X_XOR2   \PCI-PAR/$3I2493  (
    .I0(\PCI-PAR/PER_4845 ),
    .I1(\PCI-PAR/$3N2761 ),
    .O(\PCI-PAR/$3N2500 )
  );
  X_XOR4   \PCI-PAR/$2I2928  (
    .I0(\PCI-PAR/P4I ),
    .I1(\PCI-PAR/P5I ),
    .I2(\PCI-PAR/P6I ),
    .I3(\PCI-PAR/P7I ),
    .O(\PCI-PAR/PER64_4858 )
  );
  X_XOR4   \PCI-PAR/X23  (
    .I0(AD60),
    .I1(AD61),
    .I2(AD62),
    .I3(AD63),
    .O(\PCI-PAR/X15I )
  );
  X_XOR3   \PCI-PAR/X22  (
    .I0(\PCI-PAR/X14I ),
    .I1(CBE_IN7),
    .I2(\PCI-PAR/X15I ),
    .O(\PCI-PAR/P7I )
  );
  X_XOR3   \PCI-PAR/X19  (
    .I0(\PCI-PAR/X12I ),
    .I1(CBE_IN6),
    .I2(\PCI-PAR/X13I ),
    .O(\PCI-PAR/P6I )
  );
  X_XOR3   \PCI-PAR/X16  (
    .I0(\PCI-PAR/X10I ),
    .I1(CBE_IN5),
    .I2(\PCI-PAR/X11I ),
    .O(\PCI-PAR/P5I )
  );
  X_XOR3   \PCI-PAR/X13  (
    .I0(\PCI-PAR/X8I ),
    .I1(CBE_IN4),
    .I2(\PCI-PAR/X9I ),
    .O(\PCI-PAR/P4I )
  );
  X_XOR4   \PCI-PAR/X12  (
    .I0(AD32),
    .I1(AD33),
    .I2(AD34),
    .I3(AD35),
    .O(\PCI-PAR/X8I )
  );
  X_XOR4   \PCI-PAR/X14  (
    .I0(AD36),
    .I1(AD37),
    .I2(AD38),
    .I3(AD39),
    .O(\PCI-PAR/X9I )
  );
  X_XOR4   \PCI-PAR/X17  (
    .I0(AD44),
    .I1(AD45),
    .I2(AD46),
    .I3(AD47),
    .O(\PCI-PAR/X11I )
  );
  X_XOR4   \PCI-PAR/X15  (
    .I0(AD40),
    .I1(AD41),
    .I2(AD42),
    .I3(AD43),
    .O(\PCI-PAR/X10I )
  );
  X_XOR4   \PCI-PAR/X18  (
    .I0(AD48),
    .I1(AD49),
    .I2(AD50),
    .I3(AD51),
    .O(\PCI-PAR/X12I )
  );
  X_XOR4   \PCI-PAR/X20  (
    .I0(AD52),
    .I1(AD53),
    .I2(AD54),
    .I3(AD55),
    .O(\PCI-PAR/X13I )
  );
  X_XOR4   \PCI-PAR/X21  (
    .I0(AD56),
    .I1(AD57),
    .I2(AD58),
    .I3(AD59),
    .O(\PCI-PAR/X14I )
  );
  X_XOR4   \PCI-PAR/$1I2751  (
    .I0(\PCI-PAR/P0I ),
    .I1(\PCI-PAR/P1I ),
    .I2(\PCI-PAR/P2I ),
    .I3(\PCI-PAR/P3I ),
    .O(\PCI-PAR/PER_4845 )
  );
  X_XOR3   \PCI-PAR/X1  (
    .I0(\PCI-PAR/X0I ),
    .I1(CBE_IN0),
    .I2(\PCI-PAR/X1I ),
    .O(\PCI-PAR/P0I )
  );
  X_XOR4   \PCI-PAR/X0  (
    .I0(AD0),
    .I1(AD1),
    .I2(AD2),
    .I3(AD3),
    .O(\PCI-PAR/X0I )
  );
  X_XOR4   \PCI-PAR/X2  (
    .I0(AD4),
    .I1(AD5),
    .I2(AD6),
    .I3(AD7),
    .O(\PCI-PAR/X1I )
  );
  X_XOR3   \PCI-PAR/X4  (
    .I0(\PCI-PAR/X2I ),
    .I1(CBE_IN1),
    .I2(\PCI-PAR/X3I ),
    .O(\PCI-PAR/P1I )
  );
  X_XOR4   \PCI-PAR/X3  (
    .I0(AD8),
    .I1(AD9),
    .I2(AD10),
    .I3(AD11),
    .O(\PCI-PAR/X2I )
  );
  X_XOR4   \PCI-PAR/X5  (
    .I0(AD12),
    .I1(AD13),
    .I2(AD14),
    .I3(AD15),
    .O(\PCI-PAR/X3I )
  );
  X_XOR3   \PCI-PAR/X7  (
    .I0(\PCI-PAR/X4I ),
    .I1(CBE_IN2),
    .I2(\PCI-PAR/X5I ),
    .O(\PCI-PAR/P2I )
  );
  X_XOR4   \PCI-PAR/X6  (
    .I0(AD16),
    .I1(AD17),
    .I2(AD18),
    .I3(AD19),
    .O(\PCI-PAR/X4I )
  );
  X_XOR4   \PCI-PAR/X8  (
    .I0(AD20),
    .I1(AD21),
    .I2(AD22),
    .I3(AD23),
    .O(\PCI-PAR/X5I )
  );
  X_XOR3   \PCI-PAR/X10  (
    .I0(\PCI-PAR/X6I ),
    .I1(CBE_IN3),
    .I2(\PCI-PAR/X7I ),
    .O(\PCI-PAR/P3I )
  );
  X_XOR4   \PCI-PAR/X9  (
    .I0(AD24),
    .I1(AD25),
    .I2(AD26),
    .I3(AD27),
    .O(\PCI-PAR/X6I )
  );
  X_XOR4   \PCI-PAR/X11  (
    .I0(AD28),
    .I1(AD29),
    .I2(AD30),
    .I3(AD31),
    .O(\PCI-PAR/X7I )
  );
  X_ONE   \PCI-PAR/$3I3033/$1I2220  (
    .O(\PCI-PAR/$3I3033/$1N2216 )
  );
  X_BUF   \PCI-PAR/$3I3033/H  (
    .I(\PCI-PAR/$3I3033/$1N2216 ),
    .O(\PCI-PAR/$3N3020 )
  );
  X_ZERO   \PCI-PAR/$3I3034/$1I2218  (
    .O(\PCI-PAR/$3I3034/$1N2216 )
  );
  X_BUF   \PCI-PAR/$3I3034/L  (
    .I(\PCI-PAR/$3I3034/$1N2216 ),
    .O(\PCI-PAR/$3N2761 )
  );
  X_ZERO   \PCI-PAR/$4I3135/$1I2218  (
    .O(\PCI-PAR/$4I3135/$1N2216 )
  );
  X_BUF   \PCI-PAR/$4I3135/L  (
    .I(\PCI-PAR/$4I3135/$1N2216 ),
    .O(\PCI-PAR/$4N3125 )
  );
  X_ONE   \PCI-PAR/$4I3136/$1I2220  (
    .O(\PCI-PAR/$4I3136/$1N2216 )
  );
  X_BUF   \PCI-PAR/$4I3136/H  (
    .I(\PCI-PAR/$4I3136/$1N2216 ),
    .O(\PCI-PAR/$4N3107 )
  );
  X_ONE   \PCI-PAR/$7I2990/$1I2220  (
    .O(\PCI-PAR/$7I2990/$1N2216 )
  );
  X_BUF   \PCI-PAR/$7I2990/H  (
    .I(\PCI-PAR/$7I2990/$1N2216 ),
    .O(\PCI-PAR/$7N2992 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2991/UPPER/Q15  (
    .CE(\PCI-PAR/$7N2992 ),
    .CLK(CLK),
    .I(ADOUT63),
    .O(\PCI-PAR/DOQ63 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2991/UPPER/Q9  (
    .CE(\PCI-PAR/$7N2992 ),
    .CLK(CLK),
    .I(ADOUT57),
    .O(\PCI-PAR/DOQ57 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2991/UPPER/Q13  (
    .CE(\PCI-PAR/$7N2992 ),
    .CLK(CLK),
    .I(ADOUT61),
    .O(\PCI-PAR/DOQ61 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2991/UPPER/Q10  (
    .CE(\PCI-PAR/$7N2992 ),
    .CLK(CLK),
    .I(ADOUT58),
    .O(\PCI-PAR/DOQ58 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2991/UPPER/Q14  (
    .CE(\PCI-PAR/$7N2992 ),
    .CLK(CLK),
    .I(ADOUT62),
    .O(\PCI-PAR/DOQ62 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2991/UPPER/Q12  (
    .CE(\PCI-PAR/$7N2992 ),
    .CLK(CLK),
    .I(ADOUT60),
    .O(\PCI-PAR/DOQ60 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2991/UPPER/Q11  (
    .CE(\PCI-PAR/$7N2992 ),
    .CLK(CLK),
    .I(ADOUT59),
    .O(\PCI-PAR/DOQ59 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2991/UPPER/Q8  (
    .CE(\PCI-PAR/$7N2992 ),
    .CLK(CLK),
    .I(ADOUT56),
    .O(\PCI-PAR/DOQ56 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2991/UPPER/Q7  (
    .CE(\PCI-PAR/$7N2992 ),
    .CLK(CLK),
    .I(ADOUT55),
    .O(\PCI-PAR/DOQ55 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2991/UPPER/Q1  (
    .CE(\PCI-PAR/$7N2992 ),
    .CLK(CLK),
    .I(ADOUT49),
    .O(\PCI-PAR/DOQ49 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2991/UPPER/Q5  (
    .CE(\PCI-PAR/$7N2992 ),
    .CLK(CLK),
    .I(ADOUT53),
    .O(\PCI-PAR/DOQ53 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2991/UPPER/Q3  (
    .CE(\PCI-PAR/$7N2992 ),
    .CLK(CLK),
    .I(ADOUT51),
    .O(\PCI-PAR/DOQ51 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2991/UPPER/Q0  (
    .CE(\PCI-PAR/$7N2992 ),
    .CLK(CLK),
    .I(ADOUT48),
    .O(\PCI-PAR/DOQ48 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2991/UPPER/Q2  (
    .CE(\PCI-PAR/$7N2992 ),
    .CLK(CLK),
    .I(ADOUT50),
    .O(\PCI-PAR/DOQ50 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2991/UPPER/Q4  (
    .CE(\PCI-PAR/$7N2992 ),
    .CLK(CLK),
    .I(ADOUT52),
    .O(\PCI-PAR/DOQ52 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2991/UPPER/Q6  (
    .CE(\PCI-PAR/$7N2992 ),
    .CLK(CLK),
    .I(ADOUT54),
    .O(\PCI-PAR/DOQ54 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2991/LOWER/Q15  (
    .CE(\PCI-PAR/$7N2992 ),
    .CLK(CLK),
    .I(ADOUT47),
    .O(\PCI-PAR/DOQ47 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2991/LOWER/Q9  (
    .CE(\PCI-PAR/$7N2992 ),
    .CLK(CLK),
    .I(ADOUT41),
    .O(\PCI-PAR/DOQ41 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2991/LOWER/Q13  (
    .CE(\PCI-PAR/$7N2992 ),
    .CLK(CLK),
    .I(ADOUT45),
    .O(\PCI-PAR/DOQ45 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2991/LOWER/Q10  (
    .CE(\PCI-PAR/$7N2992 ),
    .CLK(CLK),
    .I(ADOUT42),
    .O(\PCI-PAR/DOQ42 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2991/LOWER/Q14  (
    .CE(\PCI-PAR/$7N2992 ),
    .CLK(CLK),
    .I(ADOUT46),
    .O(\PCI-PAR/DOQ46 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2991/LOWER/Q12  (
    .CE(\PCI-PAR/$7N2992 ),
    .CLK(CLK),
    .I(ADOUT44),
    .O(\PCI-PAR/DOQ44 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2991/LOWER/Q11  (
    .CE(\PCI-PAR/$7N2992 ),
    .CLK(CLK),
    .I(ADOUT43),
    .O(\PCI-PAR/DOQ43 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2991/LOWER/Q8  (
    .CE(\PCI-PAR/$7N2992 ),
    .CLK(CLK),
    .I(ADOUT40),
    .O(\PCI-PAR/DOQ40 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2991/LOWER/Q7  (
    .CE(\PCI-PAR/$7N2992 ),
    .CLK(CLK),
    .I(ADOUT39),
    .O(\PCI-PAR/DOQ39 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2991/LOWER/Q1  (
    .CE(\PCI-PAR/$7N2992 ),
    .CLK(CLK),
    .I(ADOUT33),
    .O(\PCI-PAR/DOQ33 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2991/LOWER/Q5  (
    .CE(\PCI-PAR/$7N2992 ),
    .CLK(CLK),
    .I(ADOUT37),
    .O(\PCI-PAR/DOQ37 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2991/LOWER/Q3  (
    .CE(\PCI-PAR/$7N2992 ),
    .CLK(CLK),
    .I(ADOUT35),
    .O(\PCI-PAR/DOQ35 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2991/LOWER/Q0  (
    .CE(\PCI-PAR/$7N2992 ),
    .CLK(CLK),
    .I(ADOUT32),
    .O(\PCI-PAR/DOQ32 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2991/LOWER/Q2  (
    .CE(\PCI-PAR/$7N2992 ),
    .CLK(CLK),
    .I(ADOUT34),
    .O(\PCI-PAR/DOQ34 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2991/LOWER/Q4  (
    .CE(\PCI-PAR/$7N2992 ),
    .CLK(CLK),
    .I(ADOUT36),
    .O(\PCI-PAR/DOQ36 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2991/LOWER/Q6  (
    .CE(\PCI-PAR/$7N2992 ),
    .CLK(CLK),
    .I(ADOUT38),
    .O(\PCI-PAR/DOQ38 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2996/UPPER/Q15  (
    .CE(\PCI-PAR/$7N2995 ),
    .CLK(CLK),
    .I(ADOUT31),
    .O(\PCI-PAR/DOQ31 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2996/UPPER/Q9  (
    .CE(\PCI-PAR/$7N2995 ),
    .CLK(CLK),
    .I(ADOUT25),
    .O(\PCI-PAR/DOQ25 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2996/UPPER/Q13  (
    .CE(\PCI-PAR/$7N2995 ),
    .CLK(CLK),
    .I(ADOUT29),
    .O(\PCI-PAR/DOQ29 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2996/UPPER/Q10  (
    .CE(\PCI-PAR/$7N2995 ),
    .CLK(CLK),
    .I(ADOUT26),
    .O(\PCI-PAR/DOQ26 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2996/UPPER/Q14  (
    .CE(\PCI-PAR/$7N2995 ),
    .CLK(CLK),
    .I(ADOUT30),
    .O(\PCI-PAR/DOQ30 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2996/UPPER/Q12  (
    .CE(\PCI-PAR/$7N2995 ),
    .CLK(CLK),
    .I(ADOUT28),
    .O(\PCI-PAR/DOQ28 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2996/UPPER/Q11  (
    .CE(\PCI-PAR/$7N2995 ),
    .CLK(CLK),
    .I(ADOUT27),
    .O(\PCI-PAR/DOQ27 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2996/UPPER/Q8  (
    .CE(\PCI-PAR/$7N2995 ),
    .CLK(CLK),
    .I(ADOUT24),
    .O(\PCI-PAR/DOQ24 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2996/UPPER/Q7  (
    .CE(\PCI-PAR/$7N2995 ),
    .CLK(CLK),
    .I(ADOUT23),
    .O(\PCI-PAR/DOQ23 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2996/UPPER/Q1  (
    .CE(\PCI-PAR/$7N2995 ),
    .CLK(CLK),
    .I(ADOUT17),
    .O(\PCI-PAR/DOQ17 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2996/UPPER/Q5  (
    .CE(\PCI-PAR/$7N2995 ),
    .CLK(CLK),
    .I(ADOUT21),
    .O(\PCI-PAR/DOQ21 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2996/UPPER/Q3  (
    .CE(\PCI-PAR/$7N2995 ),
    .CLK(CLK),
    .I(ADOUT19),
    .O(\PCI-PAR/DOQ19 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2996/UPPER/Q0  (
    .CE(\PCI-PAR/$7N2995 ),
    .CLK(CLK),
    .I(ADOUT16),
    .O(\PCI-PAR/DOQ16 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2996/UPPER/Q2  (
    .CE(\PCI-PAR/$7N2995 ),
    .CLK(CLK),
    .I(ADOUT18),
    .O(\PCI-PAR/DOQ18 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2996/UPPER/Q4  (
    .CE(\PCI-PAR/$7N2995 ),
    .CLK(CLK),
    .I(ADOUT20),
    .O(\PCI-PAR/DOQ20 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2996/UPPER/Q6  (
    .CE(\PCI-PAR/$7N2995 ),
    .CLK(CLK),
    .I(ADOUT22),
    .O(\PCI-PAR/DOQ22 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2996/LOWER/Q15  (
    .CE(\PCI-PAR/$7N2995 ),
    .CLK(CLK),
    .I(ADOUT15),
    .O(\PCI-PAR/DOQ15 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2996/LOWER/Q9  (
    .CE(\PCI-PAR/$7N2995 ),
    .CLK(CLK),
    .I(ADOUT9),
    .O(\PCI-PAR/DOQ9 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2996/LOWER/Q13  (
    .CE(\PCI-PAR/$7N2995 ),
    .CLK(CLK),
    .I(ADOUT13),
    .O(\PCI-PAR/DOQ13 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2996/LOWER/Q10  (
    .CE(\PCI-PAR/$7N2995 ),
    .CLK(CLK),
    .I(ADOUT10),
    .O(\PCI-PAR/DOQ10 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2996/LOWER/Q14  (
    .CE(\PCI-PAR/$7N2995 ),
    .CLK(CLK),
    .I(ADOUT14),
    .O(\PCI-PAR/DOQ14 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2996/LOWER/Q12  (
    .CE(\PCI-PAR/$7N2995 ),
    .CLK(CLK),
    .I(ADOUT12),
    .O(\PCI-PAR/DOQ12 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2996/LOWER/Q11  (
    .CE(\PCI-PAR/$7N2995 ),
    .CLK(CLK),
    .I(ADOUT11),
    .O(\PCI-PAR/DOQ11 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2996/LOWER/Q8  (
    .CE(\PCI-PAR/$7N2995 ),
    .CLK(CLK),
    .I(ADOUT8),
    .O(\PCI-PAR/DOQ8 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2996/LOWER/Q7  (
    .CE(\PCI-PAR/$7N2995 ),
    .CLK(CLK),
    .I(ADOUT7),
    .O(\PCI-PAR/DOQ7 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2996/LOWER/Q1  (
    .CE(\PCI-PAR/$7N2995 ),
    .CLK(CLK),
    .I(ADOUT1),
    .O(\PCI-PAR/DOQ1 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2996/LOWER/Q5  (
    .CE(\PCI-PAR/$7N2995 ),
    .CLK(CLK),
    .I(ADOUT5),
    .O(\PCI-PAR/DOQ5 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2996/LOWER/Q3  (
    .CE(\PCI-PAR/$7N2995 ),
    .CLK(CLK),
    .I(ADOUT3),
    .O(\PCI-PAR/DOQ3 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2996/LOWER/Q0  (
    .CE(\PCI-PAR/$7N2995 ),
    .CLK(CLK),
    .I(ADOUT0),
    .O(\PCI-PAR/DOQ0 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2996/LOWER/Q2  (
    .CE(\PCI-PAR/$7N2995 ),
    .CLK(CLK),
    .I(ADOUT2),
    .O(\PCI-PAR/DOQ2 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2996/LOWER/Q4  (
    .CE(\PCI-PAR/$7N2995 ),
    .CLK(CLK),
    .I(ADOUT4),
    .O(\PCI-PAR/DOQ4 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-PAR/$7I2996/LOWER/Q6  (
    .CE(\PCI-PAR/$7N2995 ),
    .CLK(CLK),
    .I(ADOUT6),
    .O(\PCI-PAR/DOQ6 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_ONE   \PCI-PAR/$7I2997/$1I2220  (
    .O(\PCI-PAR/$7I2997/$1N2216 )
  );
  X_BUF   \PCI-PAR/$7I2997/H  (
    .I(\PCI-PAR/$7I2997/$1N2216 ),
    .O(\PCI-PAR/$7N2995 )
  );
  X_ZERO   \$3I3124/$1I2218  (
    .O(\$3I3124/$1N2216 )
  );
  X_BUF   \$3I3124/L  (
    .I(\$3I3124/$1N2216 ),
    .O(BAR7)
  );
  X_ZERO   \$3I3125/$1I2218  (
    .O(\$3I3125/$1N2216 )
  );
  X_BUF   \$3I3125/L  (
    .I(\$3I3125/$1N2216 ),
    .O(BAR6)
  );
  X_ZERO   \$3I3126/$1I2218  (
    .O(\$3I3126/$1N2216 )
  );
  X_BUF   \$3I3126/L  (
    .I(\$3I3126/$1N2216 ),
    .O(BAR5)
  );
  X_ZERO   \$3I3127/$1I2218  (
    .O(\$3I3127/$1N2216 )
  );
  X_BUF   \$3I3127/L  (
    .I(\$3I3127/$1N2216 ),
    .O(BAR4)
  );
  X_ZERO   \$3I3128/$1I2218  (
    .O(\$3I3128/$1N2216 )
  );
  X_BUF   \$3I3128/L  (
    .I(\$3I3128/$1N2216 ),
    .O(BAR3)
  );
  X_ZERO   \$3I3355/$1I2218  (
    .O(\$3I3355/$1N2216 )
  );
  X_BUF   \$3I3355/L  (
    .I(\$3I3355/$1N2216 ),
    .O(NL7)
  );
  X_ZERO   \$3I3356/$1I2218  (
    .O(\$3I3356/$1N2216 )
  );
  X_BUF   \$3I3356/L  (
    .I(\$3I3356/$1N2216 ),
    .O(NL6)
  );
  X_ZERO   \$3I3357/$1I2218  (
    .O(\$3I3357/$1N2216 )
  );
  X_BUF   \$3I3357/L  (
    .I(\$3I3357/$1N2216 ),
    .O(NL5)
  );
  X_ZERO   \$3I3358/$1I2218  (
    .O(\$3I3358/$1N2216 )
  );
  X_BUF   \$3I3358/L  (
    .I(\$3I3358/$1N2216 ),
    .O(NL4)
  );
  X_ZERO   \$3I3359/$1I2218  (
    .O(\$3I3359/$1N2216 )
  );
  X_BUF   \$3I3359/L  (
    .I(\$3I3359/$1N2216 ),
    .O(NL3)
  );
  X_TRI   \4/UPPER/T0  (
    .I(\0BR16 ),
    .O(ADIO16),
    .CTL(\NlwInverterSignal_4/UPPER/T0/T )
  );
  X_TRI   \4/UPPER/T1  (
    .I(\0BR17 ),
    .O(ADIO17),
    .CTL(\NlwInverterSignal_4/UPPER/T1/T )
  );
  X_TRI   \4/UPPER/T2  (
    .I(\0BR18 ),
    .O(ADIO18),
    .CTL(\NlwInverterSignal_4/UPPER/T2/T )
  );
  X_TRI   \4/UPPER/T3  (
    .I(\0BR19 ),
    .O(ADIO19),
    .CTL(\NlwInverterSignal_4/UPPER/T3/T )
  );
  X_TRI   \4/UPPER/T4  (
    .I(\0BR20 ),
    .O(ADIO20),
    .CTL(\NlwInverterSignal_4/UPPER/T4/T )
  );
  X_TRI   \4/UPPER/T5  (
    .I(\0BR21 ),
    .O(ADIO21),
    .CTL(\NlwInverterSignal_4/UPPER/T5/T )
  );
  X_TRI   \4/UPPER/T6  (
    .I(\0BR22 ),
    .O(ADIO22),
    .CTL(\NlwInverterSignal_4/UPPER/T6/T )
  );
  X_TRI   \4/UPPER/T7  (
    .I(\0BR23 ),
    .O(ADIO23),
    .CTL(\NlwInverterSignal_4/UPPER/T7/T )
  );
  X_TRI   \4/UPPER/T8  (
    .I(\0BR24 ),
    .O(ADIO24),
    .CTL(\NlwInverterSignal_4/UPPER/T8/T )
  );
  X_TRI   \4/UPPER/T9  (
    .I(\0BR25 ),
    .O(ADIO25),
    .CTL(\NlwInverterSignal_4/UPPER/T9/T )
  );
  X_TRI   \4/UPPER/T10  (
    .I(\0BR26 ),
    .O(ADIO26),
    .CTL(\NlwInverterSignal_4/UPPER/T10/T )
  );
  X_TRI   \4/UPPER/T11  (
    .I(\0BR27 ),
    .O(ADIO27),
    .CTL(\NlwInverterSignal_4/UPPER/T11/T )
  );
  X_TRI   \4/UPPER/T12  (
    .I(\0BR28 ),
    .O(ADIO28),
    .CTL(\NlwInverterSignal_4/UPPER/T12/T )
  );
  X_TRI   \4/UPPER/T13  (
    .I(\0BR29 ),
    .O(ADIO29),
    .CTL(\NlwInverterSignal_4/UPPER/T13/T )
  );
  X_TRI   \4/UPPER/T14  (
    .I(\0BR30 ),
    .O(ADIO30),
    .CTL(\NlwInverterSignal_4/UPPER/T14/T )
  );
  X_TRI   \4/UPPER/T15  (
    .I(\0BR31 ),
    .O(ADIO31),
    .CTL(\NlwInverterSignal_4/UPPER/T15/T )
  );
  X_TRI   \4/LOWER/T0  (
    .I(\0BR0 ),
    .O(ADIO0),
    .CTL(\NlwInverterSignal_4/LOWER/T0/T )
  );
  X_TRI   \4/LOWER/T1  (
    .I(\0BR1 ),
    .O(ADIO1),
    .CTL(\NlwInverterSignal_4/LOWER/T1/T )
  );
  X_TRI   \4/LOWER/T2  (
    .I(\0BR2 ),
    .O(ADIO2),
    .CTL(\NlwInverterSignal_4/LOWER/T2/T )
  );
  X_TRI   \4/LOWER/T3  (
    .I(\0BR3 ),
    .O(ADIO3),
    .CTL(\NlwInverterSignal_4/LOWER/T3/T )
  );
  X_TRI   \4/LOWER/T4  (
    .I(\0BR4 ),
    .O(ADIO4),
    .CTL(\NlwInverterSignal_4/LOWER/T4/T )
  );
  X_TRI   \4/LOWER/T5  (
    .I(\0BR5 ),
    .O(ADIO5),
    .CTL(\NlwInverterSignal_4/LOWER/T5/T )
  );
  X_TRI   \4/LOWER/T6  (
    .I(\0BR6 ),
    .O(ADIO6),
    .CTL(\NlwInverterSignal_4/LOWER/T6/T )
  );
  X_TRI   \4/LOWER/T7  (
    .I(\0BR7 ),
    .O(ADIO7),
    .CTL(\NlwInverterSignal_4/LOWER/T7/T )
  );
  X_TRI   \4/LOWER/T8  (
    .I(\0BR8 ),
    .O(ADIO8),
    .CTL(\NlwInverterSignal_4/LOWER/T8/T )
  );
  X_TRI   \4/LOWER/T9  (
    .I(\0BR9 ),
    .O(ADIO9),
    .CTL(\NlwInverterSignal_4/LOWER/T9/T )
  );
  X_TRI   \4/LOWER/T10  (
    .I(\0BR10 ),
    .O(ADIO10),
    .CTL(\NlwInverterSignal_4/LOWER/T10/T )
  );
  X_TRI   \4/LOWER/T11  (
    .I(\0BR11 ),
    .O(ADIO11),
    .CTL(\NlwInverterSignal_4/LOWER/T11/T )
  );
  X_TRI   \4/LOWER/T12  (
    .I(\0BR12 ),
    .O(ADIO12),
    .CTL(\NlwInverterSignal_4/LOWER/T12/T )
  );
  X_TRI   \4/LOWER/T13  (
    .I(\0BR13 ),
    .O(ADIO13),
    .CTL(\NlwInverterSignal_4/LOWER/T13/T )
  );
  X_TRI   \4/LOWER/T14  (
    .I(\0BR14 ),
    .O(ADIO14),
    .CTL(\NlwInverterSignal_4/LOWER/T14/T )
  );
  X_TRI   \4/LOWER/T15  (
    .I(\0BR15 ),
    .O(ADIO15),
    .CTL(\NlwInverterSignal_4/LOWER/T15/T )
  );
  X_TRI   \5/UPPER/T0  (
    .I(\1BR16 ),
    .O(ADIO16),
    .CTL(\NlwInverterSignal_5/UPPER/T0/T )
  );
  X_TRI   \5/UPPER/T1  (
    .I(\1BR17 ),
    .O(ADIO17),
    .CTL(\NlwInverterSignal_5/UPPER/T1/T )
  );
  X_TRI   \5/UPPER/T2  (
    .I(\1BR18 ),
    .O(ADIO18),
    .CTL(\NlwInverterSignal_5/UPPER/T2/T )
  );
  X_TRI   \5/UPPER/T3  (
    .I(\1BR19 ),
    .O(ADIO19),
    .CTL(\NlwInverterSignal_5/UPPER/T3/T )
  );
  X_TRI   \5/UPPER/T4  (
    .I(\1BR20 ),
    .O(ADIO20),
    .CTL(\NlwInverterSignal_5/UPPER/T4/T )
  );
  X_TRI   \5/UPPER/T5  (
    .I(\1BR21 ),
    .O(ADIO21),
    .CTL(\NlwInverterSignal_5/UPPER/T5/T )
  );
  X_TRI   \5/UPPER/T6  (
    .I(\1BR22 ),
    .O(ADIO22),
    .CTL(\NlwInverterSignal_5/UPPER/T6/T )
  );
  X_TRI   \5/UPPER/T7  (
    .I(\1BR23 ),
    .O(ADIO23),
    .CTL(\NlwInverterSignal_5/UPPER/T7/T )
  );
  X_TRI   \5/UPPER/T8  (
    .I(\1BR24 ),
    .O(ADIO24),
    .CTL(\NlwInverterSignal_5/UPPER/T8/T )
  );
  X_TRI   \5/UPPER/T9  (
    .I(\1BR25 ),
    .O(ADIO25),
    .CTL(\NlwInverterSignal_5/UPPER/T9/T )
  );
  X_TRI   \5/UPPER/T10  (
    .I(\1BR26 ),
    .O(ADIO26),
    .CTL(\NlwInverterSignal_5/UPPER/T10/T )
  );
  X_TRI   \5/UPPER/T11  (
    .I(\1BR27 ),
    .O(ADIO27),
    .CTL(\NlwInverterSignal_5/UPPER/T11/T )
  );
  X_TRI   \5/UPPER/T12  (
    .I(\1BR28 ),
    .O(ADIO28),
    .CTL(\NlwInverterSignal_5/UPPER/T12/T )
  );
  X_TRI   \5/UPPER/T13  (
    .I(\1BR29 ),
    .O(ADIO29),
    .CTL(\NlwInverterSignal_5/UPPER/T13/T )
  );
  X_TRI   \5/UPPER/T14  (
    .I(\1BR30 ),
    .O(ADIO30),
    .CTL(\NlwInverterSignal_5/UPPER/T14/T )
  );
  X_TRI   \5/UPPER/T15  (
    .I(\1BR31 ),
    .O(ADIO31),
    .CTL(\NlwInverterSignal_5/UPPER/T15/T )
  );
  X_TRI   \5/LOWER/T0  (
    .I(\1BR0 ),
    .O(ADIO0),
    .CTL(\NlwInverterSignal_5/LOWER/T0/T )
  );
  X_TRI   \5/LOWER/T1  (
    .I(\1BR1 ),
    .O(ADIO1),
    .CTL(\NlwInverterSignal_5/LOWER/T1/T )
  );
  X_TRI   \5/LOWER/T2  (
    .I(\1BR2 ),
    .O(ADIO2),
    .CTL(\NlwInverterSignal_5/LOWER/T2/T )
  );
  X_TRI   \5/LOWER/T3  (
    .I(\1BR3 ),
    .O(ADIO3),
    .CTL(\NlwInverterSignal_5/LOWER/T3/T )
  );
  X_TRI   \5/LOWER/T4  (
    .I(\1BR4 ),
    .O(ADIO4),
    .CTL(\NlwInverterSignal_5/LOWER/T4/T )
  );
  X_TRI   \5/LOWER/T5  (
    .I(\1BR5 ),
    .O(ADIO5),
    .CTL(\NlwInverterSignal_5/LOWER/T5/T )
  );
  X_TRI   \5/LOWER/T6  (
    .I(\1BR6 ),
    .O(ADIO6),
    .CTL(\NlwInverterSignal_5/LOWER/T6/T )
  );
  X_TRI   \5/LOWER/T7  (
    .I(\1BR7 ),
    .O(ADIO7),
    .CTL(\NlwInverterSignal_5/LOWER/T7/T )
  );
  X_TRI   \5/LOWER/T8  (
    .I(\1BR8 ),
    .O(ADIO8),
    .CTL(\NlwInverterSignal_5/LOWER/T8/T )
  );
  X_TRI   \5/LOWER/T9  (
    .I(\1BR9 ),
    .O(ADIO9),
    .CTL(\NlwInverterSignal_5/LOWER/T9/T )
  );
  X_TRI   \5/LOWER/T10  (
    .I(\1BR10 ),
    .O(ADIO10),
    .CTL(\NlwInverterSignal_5/LOWER/T10/T )
  );
  X_TRI   \5/LOWER/T11  (
    .I(\1BR11 ),
    .O(ADIO11),
    .CTL(\NlwInverterSignal_5/LOWER/T11/T )
  );
  X_TRI   \5/LOWER/T12  (
    .I(\1BR12 ),
    .O(ADIO12),
    .CTL(\NlwInverterSignal_5/LOWER/T12/T )
  );
  X_TRI   \5/LOWER/T13  (
    .I(\1BR13 ),
    .O(ADIO13),
    .CTL(\NlwInverterSignal_5/LOWER/T13/T )
  );
  X_TRI   \5/LOWER/T14  (
    .I(\1BR14 ),
    .O(ADIO14),
    .CTL(\NlwInverterSignal_5/LOWER/T14/T )
  );
  X_TRI   \5/LOWER/T15  (
    .I(\1BR15 ),
    .O(ADIO15),
    .CTL(\NlwInverterSignal_5/LOWER/T15/T )
  );
  X_TRI   \6/UPPER/T0  (
    .I(\2BR16 ),
    .O(ADIO16),
    .CTL(\NlwInverterSignal_6/UPPER/T0/T )
  );
  X_TRI   \6/UPPER/T1  (
    .I(\2BR17 ),
    .O(ADIO17),
    .CTL(\NlwInverterSignal_6/UPPER/T1/T )
  );
  X_TRI   \6/UPPER/T2  (
    .I(\2BR18 ),
    .O(ADIO18),
    .CTL(\NlwInverterSignal_6/UPPER/T2/T )
  );
  X_TRI   \6/UPPER/T3  (
    .I(\2BR19 ),
    .O(ADIO19),
    .CTL(\NlwInverterSignal_6/UPPER/T3/T )
  );
  X_TRI   \6/UPPER/T4  (
    .I(\2BR20 ),
    .O(ADIO20),
    .CTL(\NlwInverterSignal_6/UPPER/T4/T )
  );
  X_TRI   \6/UPPER/T5  (
    .I(\2BR21 ),
    .O(ADIO21),
    .CTL(\NlwInverterSignal_6/UPPER/T5/T )
  );
  X_TRI   \6/UPPER/T6  (
    .I(\2BR22 ),
    .O(ADIO22),
    .CTL(\NlwInverterSignal_6/UPPER/T6/T )
  );
  X_TRI   \6/UPPER/T7  (
    .I(\2BR23 ),
    .O(ADIO23),
    .CTL(\NlwInverterSignal_6/UPPER/T7/T )
  );
  X_TRI   \6/UPPER/T8  (
    .I(\2BR24 ),
    .O(ADIO24),
    .CTL(\NlwInverterSignal_6/UPPER/T8/T )
  );
  X_TRI   \6/UPPER/T9  (
    .I(\2BR25 ),
    .O(ADIO25),
    .CTL(\NlwInverterSignal_6/UPPER/T9/T )
  );
  X_TRI   \6/UPPER/T10  (
    .I(\2BR26 ),
    .O(ADIO26),
    .CTL(\NlwInverterSignal_6/UPPER/T10/T )
  );
  X_TRI   \6/UPPER/T11  (
    .I(\2BR27 ),
    .O(ADIO27),
    .CTL(\NlwInverterSignal_6/UPPER/T11/T )
  );
  X_TRI   \6/UPPER/T12  (
    .I(\2BR28 ),
    .O(ADIO28),
    .CTL(\NlwInverterSignal_6/UPPER/T12/T )
  );
  X_TRI   \6/UPPER/T13  (
    .I(\2BR29 ),
    .O(ADIO29),
    .CTL(\NlwInverterSignal_6/UPPER/T13/T )
  );
  X_TRI   \6/UPPER/T14  (
    .I(\2BR30 ),
    .O(ADIO30),
    .CTL(\NlwInverterSignal_6/UPPER/T14/T )
  );
  X_TRI   \6/UPPER/T15  (
    .I(\2BR31 ),
    .O(ADIO31),
    .CTL(\NlwInverterSignal_6/UPPER/T15/T )
  );
  X_TRI   \6/LOWER/T0  (
    .I(\2BR0 ),
    .O(ADIO0),
    .CTL(\NlwInverterSignal_6/LOWER/T0/T )
  );
  X_TRI   \6/LOWER/T1  (
    .I(\2BR1 ),
    .O(ADIO1),
    .CTL(\NlwInverterSignal_6/LOWER/T1/T )
  );
  X_TRI   \6/LOWER/T2  (
    .I(\2BR2 ),
    .O(ADIO2),
    .CTL(\NlwInverterSignal_6/LOWER/T2/T )
  );
  X_TRI   \6/LOWER/T3  (
    .I(\2BR3 ),
    .O(ADIO3),
    .CTL(\NlwInverterSignal_6/LOWER/T3/T )
  );
  X_TRI   \6/LOWER/T4  (
    .I(\2BR4 ),
    .O(ADIO4),
    .CTL(\NlwInverterSignal_6/LOWER/T4/T )
  );
  X_TRI   \6/LOWER/T5  (
    .I(\2BR5 ),
    .O(ADIO5),
    .CTL(\NlwInverterSignal_6/LOWER/T5/T )
  );
  X_TRI   \6/LOWER/T6  (
    .I(\2BR6 ),
    .O(ADIO6),
    .CTL(\NlwInverterSignal_6/LOWER/T6/T )
  );
  X_TRI   \6/LOWER/T7  (
    .I(\2BR7 ),
    .O(ADIO7),
    .CTL(\NlwInverterSignal_6/LOWER/T7/T )
  );
  X_TRI   \6/LOWER/T8  (
    .I(\2BR8 ),
    .O(ADIO8),
    .CTL(\NlwInverterSignal_6/LOWER/T8/T )
  );
  X_TRI   \6/LOWER/T9  (
    .I(\2BR9 ),
    .O(ADIO9),
    .CTL(\NlwInverterSignal_6/LOWER/T9/T )
  );
  X_TRI   \6/LOWER/T10  (
    .I(\2BR10 ),
    .O(ADIO10),
    .CTL(\NlwInverterSignal_6/LOWER/T10/T )
  );
  X_TRI   \6/LOWER/T11  (
    .I(\2BR11 ),
    .O(ADIO11),
    .CTL(\NlwInverterSignal_6/LOWER/T11/T )
  );
  X_TRI   \6/LOWER/T12  (
    .I(\2BR12 ),
    .O(ADIO12),
    .CTL(\NlwInverterSignal_6/LOWER/T12/T )
  );
  X_TRI   \6/LOWER/T13  (
    .I(\2BR13 ),
    .O(ADIO13),
    .CTL(\NlwInverterSignal_6/LOWER/T13/T )
  );
  X_TRI   \6/LOWER/T14  (
    .I(\2BR14 ),
    .O(ADIO14),
    .CTL(\NlwInverterSignal_6/LOWER/T14/T )
  );
  X_TRI   \6/LOWER/T15  (
    .I(\2BR15 ),
    .O(ADIO15),
    .CTL(\NlwInverterSignal_6/LOWER/T15/T )
  );
  X_BUF   \$3I3818/NC  (
    .I(NlwRenamedSig_OI_BASE_HIT7),
    .O(\NLW_$3I3818/NC_O_UNCONNECTED )
  );
  X_BUF   \$3I3819/NC  (
    .I(NlwRenamedSig_OI_BASE_HIT6),
    .O(\NLW_$3I3819/NC_O_UNCONNECTED )
  );
  X_BUF   \$3I3820/NC  (
    .I(NlwRenamedSig_OI_BASE_HIT5),
    .O(\NLW_$3I3820/NC_O_UNCONNECTED )
  );
  X_BUF   \$3I3821/NC  (
    .I(NlwRenamedSig_OI_BASE_HIT4),
    .O(\NLW_$3I3821/NC_O_UNCONNECTED )
  );
  X_BUF   \$3I3822/NC  (
    .I(NlwRenamedSig_OI_BASE_HIT3),
    .O(\NLW_$3I3822/NC_O_UNCONNECTED )
  );
  X_BUF   \$3I3823/NC  (
    .I(NlwRenamedSig_OI_BASE_HIT2),
    .O(\NLW_$3I3823/NC_O_UNCONNECTED )
  );
  X_BUF   \$3I3824/NC  (
    .I(NlwRenamedSig_OI_BASE_HIT1),
    .O(\NLW_$3I3824/NC_O_UNCONNECTED )
  );
  X_BUF   \$3I3825/NC  (
    .I(NlwRenamedSig_OI_BASE_HIT0),
    .O(\NLW_$3I3825/NC_O_UNCONNECTED )
  );
  X_BUF   \$3I3826/NC  (
    .I(NL_MEM7),
    .O(\NLW_$3I3826/NC_O_UNCONNECTED )
  );
  X_BUF   \$3I3827/NC  (
    .I(NL_MEM6),
    .O(\NLW_$3I3827/NC_O_UNCONNECTED )
  );
  X_BUF   \$3I3828/NC  (
    .I(NL_MEM5),
    .O(\NLW_$3I3828/NC_O_UNCONNECTED )
  );
  X_BUF   \$3I3829/NC  (
    .I(NL_MEM4),
    .O(\NLW_$3I3829/NC_O_UNCONNECTED )
  );
  X_BUF   \$3I3830/NC  (
    .I(NL_MEM3),
    .O(\NLW_$3I3830/NC_O_UNCONNECTED )
  );
  X_BUF   \$3I3831/NC  (
    .I(NL_MEM2),
    .O(\NLW_$3I3831/NC_O_UNCONNECTED )
  );
  X_BUF   \$3I3832/NC  (
    .I(NL_MEM1),
    .O(\NLW_$3I3832/NC_O_UNCONNECTED )
  );
  X_BUF   \$3I3833/NC  (
    .I(NL_MEM0),
    .O(\NLW_$3I3833/NC_O_UNCONNECTED )
  );
  X_AND4   \BAR0/$2I3324  (
    .I0(\BAR0/CSRENNL ),
    .I1(\BAR0/MATCH ),
    .I2(ADDR_VLD1),
    .I3(\BAR0/ENABLENL ),
    .O(\BAR0/NS_HITNL )
  );
  X_INV   \BAR0/$2I3284  (
    .I(CFG36),
    .O(\BAR0/NL_CE )
  );
  X_AND2   \BAR0/$2I3275  (
    .I0(\TSTOP_I- ),
    .I1(\BAR0/$2N3280 ),
    .O(\BAR0/NS_NL_MEM )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR0/NL  (
    .CE(\BAR0/NL_CE ),
    .CLK(CLK),
    .I(\BAR0/NS_NL_MEM ),
    .O(NL_MEM0),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_OR2   \BAR0/$2I3268  (
    .I0(\BAR0/$2N3273 ),
    .I1(NL_MEM0),
    .O(\BAR0/$2N3280 )
  );
  X_AND2   \BAR0/$2I3267  (
    .I0(\BAR0/UNALIGN ),
    .I1(\BAR0/NS_HITNL ),
    .O(\BAR0/$2N3273 )
  );
  X_OR2   \BAR0/$2I3263  (
    .I0(AD1),
    .I1(AD0),
    .O(\BAR0/UNALIGN )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR0/EQ64  (
    .CE(VCC),
    .CLK(CLK),
    .I(NS_BH64_0),
    .O(BH64_0),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR0/EQ32  (
    .CE(VCC),
    .CLK(CLK),
    .I(NS_BASE_HIT0),
    .O(NlwRenamedSig_OI_BASE_HIT0),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND4   \BAR0/$1I3455  (
    .I0(\BAR0/CSREN64 ),
    .I1(\BAR0/MATCH ),
    .I2(ADDR_VLD64),
    .I3(CFG241),
    .O(NS_BH64_0)
  );
  X_AND4   \BAR0/$1I3437  (
    .I0(\BAR0/CSREN32 ),
    .I1(\BAR0/MATCH ),
    .I2(ADDR_VLD1),
    .I3(\BAR0/ENABLE32 ),
    .O(NS_BASE_HIT0)
  );
  X_MUX2   \BAR0/BR-31-24/$1I3094  (
    .IB(\BAR0/$1N3369 ),
    .IA(\BAR0/BR-31-24/$1N3110 ),
    .O(\BAR0/BR-31-24/$1N3099 ),
    .SEL(\BAR0/BR-31-24/EQ10_5479 )
  );
  X_MUX2   \BAR0/BR-31-24/$1I3093  (
    .IB(\BAR0/BR-31-24/$1N3099 ),
    .IA(\BAR0/BR-31-24/$1N3111 ),
    .O(\BAR0/BR-31-24/$1N2993 ),
    .SEL(\BAR0/BR-31-24/EQ32_5482 )
  );
  X_XOR2   \BAR0/BR-31-24/X1  (
    .I0(\BAR0/BR-31-24/IN1 ),
    .I1(\0BR25 ),
    .O(\NlwInverterSignal_BAR0/BR-31-24/X1/O )
  );
  X_XOR2   \BAR0/BR-31-24/X3  (
    .I0(\BAR0/BR-31-24/IN3 ),
    .I1(\0BR27 ),
    .O(\NlwInverterSignal_BAR0/BR-31-24/X3/O )
  );
  X_AND2   \BAR0/BR-31-24/$1I3014  (
    .I0(CFG27),
    .I1(\BAR0/BR-31-24/RAWQ2 ),
    .O(\0BR26 )
  );
  X_AND2   \BAR0/BR-31-24/$1I3013  (
    .I0(AD26),
    .I1(CFG27),
    .O(\BAR0/BR-31-24/IN2 )
  );
  X_AND2   \BAR0/BR-31-24/$1I3012  (
    .I0(AD25),
    .I1(CFG26),
    .O(\BAR0/BR-31-24/IN1 )
  );
  X_AND2   \BAR0/BR-31-24/$1I3011  (
    .I0(CFG26),
    .I1(\BAR0/BR-31-24/RAWQ1 ),
    .O(\0BR25 )
  );
  X_AND2   \BAR0/BR-31-24/$1I3010  (
    .I0(CFG25),
    .I1(\BAR0/BR-31-24/RAWQ0 ),
    .O(\0BR24 )
  );
  X_AND2   \BAR0/BR-31-24/$1I3009  (
    .I0(CFG28),
    .I1(\BAR0/BR-31-24/RAWQ3 ),
    .O(\0BR27 )
  );
  X_AND2   \BAR0/BR-31-24/$1I3008  (
    .I0(AD27),
    .I1(CFG28),
    .O(\BAR0/BR-31-24/IN3 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR0/BR-31-24/Q3  (
    .CE(CE4_3),
    .CLK(CLK),
    .I(AD27),
    .O(\BAR0/BR-31-24/RAWQ3 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR0/BR-31-24/Q2  (
    .CE(CE4_3),
    .CLK(CLK),
    .I(AD26),
    .O(\BAR0/BR-31-24/RAWQ2 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR0/BR-31-24/Q1  (
    .CE(CE4_3),
    .CLK(CLK),
    .I(AD25),
    .O(\BAR0/BR-31-24/RAWQ1 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR0/BR-31-24/Q0  (
    .CE(CE4_3),
    .CLK(CLK),
    .I(AD24),
    .O(\BAR0/BR-31-24/RAWQ0 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \BAR0/BR-31-24/X2  (
    .I0(\BAR0/BR-31-24/IN2 ),
    .I1(\0BR26 ),
    .O(\NlwInverterSignal_BAR0/BR-31-24/X2/O )
  );
  X_XOR2   \BAR0/BR-31-24/X0  (
    .I0(\BAR0/BR-31-24/IN0 ),
    .I1(\0BR24 ),
    .O(\NlwInverterSignal_BAR0/BR-31-24/X0/O )
  );
  X_AND2   \BAR0/BR-31-24/A1  (
    .I0(\BAR0/BR-31-24/EQ2 ),
    .I1(\BAR0/BR-31-24/EQ3 ),
    .O(\BAR0/BR-31-24/EQ32_5482 )
  );
  X_AND2   \BAR0/BR-31-24/A0  (
    .I0(\BAR0/BR-31-24/EQ0 ),
    .I1(\BAR0/BR-31-24/EQ1 ),
    .O(\BAR0/BR-31-24/EQ10_5479 )
  );
  X_AND2   \BAR0/BR-31-24/$1I2999  (
    .I0(AD24),
    .I1(CFG25),
    .O(\BAR0/BR-31-24/IN0 )
  );
  X_AND2   \BAR0/BR-31-24/$1I2989  (
    .I0(AD28),
    .I1(CFG29),
    .O(\BAR0/BR-31-24/IN4 )
  );
  X_AND2   \BAR0/BR-31-24/A2  (
    .I0(\BAR0/BR-31-24/EQ4 ),
    .I1(\BAR0/BR-31-24/EQ5 ),
    .O(\BAR0/BR-31-24/EQ54_5469 )
  );
  X_MUX2   \BAR0/BR-31-24/$1I2986  (
    .IB(\BAR0/BR-31-24/$1N2992 ),
    .IA(\BAR0/BR-31-24/$1N2910 ),
    .O(\BAR0/$1N3380 ),
    .SEL(\BAR0/BR-31-24/EQ76_5472 )
  );
  X_MUX2   \BAR0/BR-31-24/$1I2985  (
    .IB(\BAR0/BR-31-24/$1N2993 ),
    .IA(\BAR0/BR-31-24/$1N2911 ),
    .O(\BAR0/BR-31-24/$1N2992 ),
    .SEL(\BAR0/BR-31-24/EQ54_5469 )
  );
  X_AND2   \BAR0/BR-31-24/A3  (
    .I0(\BAR0/BR-31-24/EQ6 ),
    .I1(\BAR0/BR-31-24/EQ7 ),
    .O(\BAR0/BR-31-24/EQ76_5472 )
  );
  X_XOR2   \BAR0/BR-31-24/X4  (
    .I0(\BAR0/BR-31-24/IN4 ),
    .I1(\0BR28 ),
    .O(\NlwInverterSignal_BAR0/BR-31-24/X4/O )
  );
  X_XOR2   \BAR0/BR-31-24/X6  (
    .I0(\BAR0/BR-31-24/IN6 ),
    .I1(\0BR30 ),
    .O(\NlwInverterSignal_BAR0/BR-31-24/X6/O )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR0/BR-31-24/Q4  (
    .CE(CE4_3),
    .CLK(CLK),
    .I(AD28),
    .O(\BAR0/BR-31-24/RAWQ4 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR0/BR-31-24/Q5  (
    .CE(CE4_3),
    .CLK(CLK),
    .I(AD29),
    .O(\BAR0/BR-31-24/RAWQ5 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR0/BR-31-24/Q6  (
    .CE(CE4_3),
    .CLK(CLK),
    .I(AD30),
    .O(\BAR0/BR-31-24/RAWQ6 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR0/BR-31-24/Q7  (
    .CE(CE4_3),
    .CLK(CLK),
    .I(AD31),
    .O(\BAR0/BR-31-24/RAWQ7 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND2   \BAR0/BR-31-24/$1I2960  (
    .I0(AD31),
    .I1(CFG32),
    .O(\BAR0/BR-31-24/IN7 )
  );
  X_AND2   \BAR0/BR-31-24/$1I2959  (
    .I0(CFG32),
    .I1(\BAR0/BR-31-24/RAWQ7 ),
    .O(\0BR31 )
  );
  X_AND2   \BAR0/BR-31-24/$1I2958  (
    .I0(CFG29),
    .I1(\BAR0/BR-31-24/RAWQ4 ),
    .O(\0BR28 )
  );
  X_AND2   \BAR0/BR-31-24/$1I2957  (
    .I0(CFG30),
    .I1(\BAR0/BR-31-24/RAWQ5 ),
    .O(\0BR29 )
  );
  X_AND2   \BAR0/BR-31-24/$1I2956  (
    .I0(AD29),
    .I1(CFG30),
    .O(\BAR0/BR-31-24/IN5 )
  );
  X_AND2   \BAR0/BR-31-24/$1I2955  (
    .I0(AD30),
    .I1(CFG31),
    .O(\BAR0/BR-31-24/IN6 )
  );
  X_AND2   \BAR0/BR-31-24/$1I2954  (
    .I0(CFG31),
    .I1(\BAR0/BR-31-24/RAWQ6 ),
    .O(\0BR30 )
  );
  X_XOR2   \BAR0/BR-31-24/X7  (
    .I0(\BAR0/BR-31-24/IN7 ),
    .I1(\0BR31 ),
    .O(\NlwInverterSignal_BAR0/BR-31-24/X7/O )
  );
  X_XOR2   \BAR0/BR-31-24/X5  (
    .I0(\BAR0/BR-31-24/IN5 ),
    .I1(\0BR29 ),
    .O(\NlwInverterSignal_BAR0/BR-31-24/X5/O )
  );
  X_ZERO   \BAR0/BR-31-24/$1I2909/$1I2218  (
    .O(\BAR0/BR-31-24/$1I2909/$1N2216 )
  );
  X_BUF   \BAR0/BR-31-24/$1I2909/L  (
    .I(\BAR0/BR-31-24/$1I2909/$1N2216 ),
    .O(\BAR0/BR-31-24/$1N2910 )
  );
  X_ZERO   \BAR0/BR-31-24/$1I2990/$1I2218  (
    .O(\BAR0/BR-31-24/$1I2990/$1N2216 )
  );
  X_BUF   \BAR0/BR-31-24/$1I2990/L  (
    .I(\BAR0/BR-31-24/$1I2990/$1N2216 ),
    .O(\BAR0/BR-31-24/$1N2911 )
  );
  X_ZERO   \BAR0/BR-31-24/$1I3091/$1I2218  (
    .O(\BAR0/BR-31-24/$1I3091/$1N2216 )
  );
  X_BUF   \BAR0/BR-31-24/$1I3091/L  (
    .I(\BAR0/BR-31-24/$1I3091/$1N2216 ),
    .O(\BAR0/BR-31-24/$1N3110 )
  );
  X_ZERO   \BAR0/BR-31-24/$1I3096/$1I2218  (
    .O(\BAR0/BR-31-24/$1I3096/$1N2216 )
  );
  X_BUF   \BAR0/BR-31-24/$1I3096/L  (
    .I(\BAR0/BR-31-24/$1I3096/$1N2216 ),
    .O(\BAR0/BR-31-24/$1N3111 )
  );
  X_MUX2   \BAR0/BR-23-16/$1I3094  (
    .IB(\BAR0/$1N3368 ),
    .IA(\BAR0/BR-23-16/$1N3110 ),
    .O(\BAR0/BR-23-16/$1N3099 ),
    .SEL(\BAR0/BR-23-16/EQ10_5551 )
  );
  X_MUX2   \BAR0/BR-23-16/$1I3093  (
    .IB(\BAR0/BR-23-16/$1N3099 ),
    .IA(\BAR0/BR-23-16/$1N3111 ),
    .O(\BAR0/BR-23-16/$1N2993 ),
    .SEL(\BAR0/BR-23-16/EQ32_5554 )
  );
  X_XOR2   \BAR0/BR-23-16/X1  (
    .I0(\BAR0/BR-23-16/IN1 ),
    .I1(\0BR17 ),
    .O(\NlwInverterSignal_BAR0/BR-23-16/X1/O )
  );
  X_XOR2   \BAR0/BR-23-16/X3  (
    .I0(\BAR0/BR-23-16/IN3 ),
    .I1(\0BR19 ),
    .O(\NlwInverterSignal_BAR0/BR-23-16/X3/O )
  );
  X_AND2   \BAR0/BR-23-16/$1I3014  (
    .I0(CFG19),
    .I1(\BAR0/BR-23-16/RAWQ2 ),
    .O(\0BR18 )
  );
  X_AND2   \BAR0/BR-23-16/$1I3013  (
    .I0(AD18),
    .I1(CFG19),
    .O(\BAR0/BR-23-16/IN2 )
  );
  X_AND2   \BAR0/BR-23-16/$1I3012  (
    .I0(AD17),
    .I1(CFG18),
    .O(\BAR0/BR-23-16/IN1 )
  );
  X_AND2   \BAR0/BR-23-16/$1I3011  (
    .I0(CFG18),
    .I1(\BAR0/BR-23-16/RAWQ1 ),
    .O(\0BR17 )
  );
  X_AND2   \BAR0/BR-23-16/$1I3010  (
    .I0(CFG17),
    .I1(\BAR0/BR-23-16/RAWQ0 ),
    .O(\0BR16 )
  );
  X_AND2   \BAR0/BR-23-16/$1I3009  (
    .I0(CFG20),
    .I1(\BAR0/BR-23-16/RAWQ3 ),
    .O(\0BR19 )
  );
  X_AND2   \BAR0/BR-23-16/$1I3008  (
    .I0(AD19),
    .I1(CFG20),
    .O(\BAR0/BR-23-16/IN3 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR0/BR-23-16/Q3  (
    .CE(CE4_2),
    .CLK(CLK),
    .I(AD19),
    .O(\BAR0/BR-23-16/RAWQ3 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR0/BR-23-16/Q2  (
    .CE(CE4_2),
    .CLK(CLK),
    .I(AD18),
    .O(\BAR0/BR-23-16/RAWQ2 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR0/BR-23-16/Q1  (
    .CE(CE4_2),
    .CLK(CLK),
    .I(AD17),
    .O(\BAR0/BR-23-16/RAWQ1 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR0/BR-23-16/Q0  (
    .CE(CE4_2),
    .CLK(CLK),
    .I(AD16),
    .O(\BAR0/BR-23-16/RAWQ0 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \BAR0/BR-23-16/X2  (
    .I0(\BAR0/BR-23-16/IN2 ),
    .I1(\0BR18 ),
    .O(\NlwInverterSignal_BAR0/BR-23-16/X2/O )
  );
  X_XOR2   \BAR0/BR-23-16/X0  (
    .I0(\BAR0/BR-23-16/IN0 ),
    .I1(\0BR16 ),
    .O(\NlwInverterSignal_BAR0/BR-23-16/X0/O )
  );
  X_AND2   \BAR0/BR-23-16/A1  (
    .I0(\BAR0/BR-23-16/EQ2 ),
    .I1(\BAR0/BR-23-16/EQ3 ),
    .O(\BAR0/BR-23-16/EQ32_5554 )
  );
  X_AND2   \BAR0/BR-23-16/A0  (
    .I0(\BAR0/BR-23-16/EQ0 ),
    .I1(\BAR0/BR-23-16/EQ1 ),
    .O(\BAR0/BR-23-16/EQ10_5551 )
  );
  X_AND2   \BAR0/BR-23-16/$1I2999  (
    .I0(AD16),
    .I1(CFG17),
    .O(\BAR0/BR-23-16/IN0 )
  );
  X_AND2   \BAR0/BR-23-16/$1I2989  (
    .I0(AD20),
    .I1(CFG21),
    .O(\BAR0/BR-23-16/IN4 )
  );
  X_AND2   \BAR0/BR-23-16/A2  (
    .I0(\BAR0/BR-23-16/EQ4 ),
    .I1(\BAR0/BR-23-16/EQ5 ),
    .O(\BAR0/BR-23-16/EQ54_5541 )
  );
  X_MUX2   \BAR0/BR-23-16/$1I2986  (
    .IB(\BAR0/BR-23-16/$1N2992 ),
    .IA(\BAR0/BR-23-16/$1N2910 ),
    .O(\BAR0/$1N3369 ),
    .SEL(\BAR0/BR-23-16/EQ76_5544 )
  );
  X_MUX2   \BAR0/BR-23-16/$1I2985  (
    .IB(\BAR0/BR-23-16/$1N2993 ),
    .IA(\BAR0/BR-23-16/$1N2911 ),
    .O(\BAR0/BR-23-16/$1N2992 ),
    .SEL(\BAR0/BR-23-16/EQ54_5541 )
  );
  X_AND2   \BAR0/BR-23-16/A3  (
    .I0(\BAR0/BR-23-16/EQ6 ),
    .I1(\BAR0/BR-23-16/EQ7 ),
    .O(\BAR0/BR-23-16/EQ76_5544 )
  );
  X_XOR2   \BAR0/BR-23-16/X4  (
    .I0(\BAR0/BR-23-16/IN4 ),
    .I1(\0BR20 ),
    .O(\NlwInverterSignal_BAR0/BR-23-16/X4/O )
  );
  X_XOR2   \BAR0/BR-23-16/X6  (
    .I0(\BAR0/BR-23-16/IN6 ),
    .I1(\0BR22 ),
    .O(\NlwInverterSignal_BAR0/BR-23-16/X6/O )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR0/BR-23-16/Q4  (
    .CE(CE4_2),
    .CLK(CLK),
    .I(AD20),
    .O(\BAR0/BR-23-16/RAWQ4 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR0/BR-23-16/Q5  (
    .CE(CE4_2),
    .CLK(CLK),
    .I(AD21),
    .O(\BAR0/BR-23-16/RAWQ5 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR0/BR-23-16/Q6  (
    .CE(CE4_2),
    .CLK(CLK),
    .I(AD22),
    .O(\BAR0/BR-23-16/RAWQ6 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR0/BR-23-16/Q7  (
    .CE(CE4_2),
    .CLK(CLK),
    .I(AD23),
    .O(\BAR0/BR-23-16/RAWQ7 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND2   \BAR0/BR-23-16/$1I2960  (
    .I0(AD23),
    .I1(CFG24),
    .O(\BAR0/BR-23-16/IN7 )
  );
  X_AND2   \BAR0/BR-23-16/$1I2959  (
    .I0(CFG24),
    .I1(\BAR0/BR-23-16/RAWQ7 ),
    .O(\0BR23 )
  );
  X_AND2   \BAR0/BR-23-16/$1I2958  (
    .I0(CFG21),
    .I1(\BAR0/BR-23-16/RAWQ4 ),
    .O(\0BR20 )
  );
  X_AND2   \BAR0/BR-23-16/$1I2957  (
    .I0(CFG22),
    .I1(\BAR0/BR-23-16/RAWQ5 ),
    .O(\0BR21 )
  );
  X_AND2   \BAR0/BR-23-16/$1I2956  (
    .I0(AD21),
    .I1(CFG22),
    .O(\BAR0/BR-23-16/IN5 )
  );
  X_AND2   \BAR0/BR-23-16/$1I2955  (
    .I0(AD22),
    .I1(CFG23),
    .O(\BAR0/BR-23-16/IN6 )
  );
  X_AND2   \BAR0/BR-23-16/$1I2954  (
    .I0(CFG23),
    .I1(\BAR0/BR-23-16/RAWQ6 ),
    .O(\0BR22 )
  );
  X_XOR2   \BAR0/BR-23-16/X7  (
    .I0(\BAR0/BR-23-16/IN7 ),
    .I1(\0BR23 ),
    .O(\NlwInverterSignal_BAR0/BR-23-16/X7/O )
  );
  X_XOR2   \BAR0/BR-23-16/X5  (
    .I0(\BAR0/BR-23-16/IN5 ),
    .I1(\0BR21 ),
    .O(\NlwInverterSignal_BAR0/BR-23-16/X5/O )
  );
  X_ZERO   \BAR0/BR-23-16/$1I2909/$1I2218  (
    .O(\BAR0/BR-23-16/$1I2909/$1N2216 )
  );
  X_BUF   \BAR0/BR-23-16/$1I2909/L  (
    .I(\BAR0/BR-23-16/$1I2909/$1N2216 ),
    .O(\BAR0/BR-23-16/$1N2910 )
  );
  X_ZERO   \BAR0/BR-23-16/$1I2990/$1I2218  (
    .O(\BAR0/BR-23-16/$1I2990/$1N2216 )
  );
  X_BUF   \BAR0/BR-23-16/$1I2990/L  (
    .I(\BAR0/BR-23-16/$1I2990/$1N2216 ),
    .O(\BAR0/BR-23-16/$1N2911 )
  );
  X_ZERO   \BAR0/BR-23-16/$1I3091/$1I2218  (
    .O(\BAR0/BR-23-16/$1I3091/$1N2216 )
  );
  X_BUF   \BAR0/BR-23-16/$1I3091/L  (
    .I(\BAR0/BR-23-16/$1I3091/$1N2216 ),
    .O(\BAR0/BR-23-16/$1N3110 )
  );
  X_ZERO   \BAR0/BR-23-16/$1I3096/$1I2218  (
    .O(\BAR0/BR-23-16/$1I3096/$1N2216 )
  );
  X_BUF   \BAR0/BR-23-16/$1I3096/L  (
    .I(\BAR0/BR-23-16/$1I3096/$1N2216 ),
    .O(\BAR0/BR-23-16/$1N3111 )
  );
  X_MUX2   \BAR0/BR-15-8/$1I3094  (
    .IB(\BAR0/$1N3366 ),
    .IA(\BAR0/BR-15-8/$1N3110 ),
    .O(\BAR0/BR-15-8/$1N3099 ),
    .SEL(\BAR0/BR-15-8/EQ10_5623 )
  );
  X_MUX2   \BAR0/BR-15-8/$1I3093  (
    .IB(\BAR0/BR-15-8/$1N3099 ),
    .IA(\BAR0/BR-15-8/$1N3111 ),
    .O(\BAR0/BR-15-8/$1N2993 ),
    .SEL(\BAR0/BR-15-8/EQ32_5626 )
  );
  X_XOR2   \BAR0/BR-15-8/X1  (
    .I0(\BAR0/BR-15-8/IN1 ),
    .I1(\0BR9 ),
    .O(\NlwInverterSignal_BAR0/BR-15-8/X1/O )
  );
  X_XOR2   \BAR0/BR-15-8/X3  (
    .I0(\BAR0/BR-15-8/IN3 ),
    .I1(\0BR11 ),
    .O(\NlwInverterSignal_BAR0/BR-15-8/X3/O )
  );
  X_AND2   \BAR0/BR-15-8/$1I3014  (
    .I0(CFG11),
    .I1(\BAR0/BR-15-8/RAWQ2 ),
    .O(\0BR10 )
  );
  X_AND2   \BAR0/BR-15-8/$1I3013  (
    .I0(AD10),
    .I1(CFG11),
    .O(\BAR0/BR-15-8/IN2 )
  );
  X_AND2   \BAR0/BR-15-8/$1I3012  (
    .I0(AD9),
    .I1(CFG10),
    .O(\BAR0/BR-15-8/IN1 )
  );
  X_AND2   \BAR0/BR-15-8/$1I3011  (
    .I0(CFG10),
    .I1(\BAR0/BR-15-8/RAWQ1 ),
    .O(\0BR9 )
  );
  X_AND2   \BAR0/BR-15-8/$1I3010  (
    .I0(CFG9),
    .I1(\BAR0/BR-15-8/RAWQ0 ),
    .O(\0BR8 )
  );
  X_AND2   \BAR0/BR-15-8/$1I3009  (
    .I0(CFG12),
    .I1(\BAR0/BR-15-8/RAWQ3 ),
    .O(\0BR11 )
  );
  X_AND2   \BAR0/BR-15-8/$1I3008  (
    .I0(AD11),
    .I1(CFG12),
    .O(\BAR0/BR-15-8/IN3 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR0/BR-15-8/Q3  (
    .CE(CE4_1),
    .CLK(CLK),
    .I(AD11),
    .O(\BAR0/BR-15-8/RAWQ3 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR0/BR-15-8/Q2  (
    .CE(CE4_1),
    .CLK(CLK),
    .I(AD10),
    .O(\BAR0/BR-15-8/RAWQ2 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR0/BR-15-8/Q1  (
    .CE(CE4_1),
    .CLK(CLK),
    .I(AD9),
    .O(\BAR0/BR-15-8/RAWQ1 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR0/BR-15-8/Q0  (
    .CE(CE4_1),
    .CLK(CLK),
    .I(AD8),
    .O(\BAR0/BR-15-8/RAWQ0 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \BAR0/BR-15-8/X2  (
    .I0(\BAR0/BR-15-8/IN2 ),
    .I1(\0BR10 ),
    .O(\NlwInverterSignal_BAR0/BR-15-8/X2/O )
  );
  X_XOR2   \BAR0/BR-15-8/X0  (
    .I0(\BAR0/BR-15-8/IN0 ),
    .I1(\0BR8 ),
    .O(\NlwInverterSignal_BAR0/BR-15-8/X0/O )
  );
  X_AND2   \BAR0/BR-15-8/A1  (
    .I0(\BAR0/BR-15-8/EQ2 ),
    .I1(\BAR0/BR-15-8/EQ3 ),
    .O(\BAR0/BR-15-8/EQ32_5626 )
  );
  X_AND2   \BAR0/BR-15-8/A0  (
    .I0(\BAR0/BR-15-8/EQ0 ),
    .I1(\BAR0/BR-15-8/EQ1 ),
    .O(\BAR0/BR-15-8/EQ10_5623 )
  );
  X_AND2   \BAR0/BR-15-8/$1I2999  (
    .I0(AD8),
    .I1(CFG9),
    .O(\BAR0/BR-15-8/IN0 )
  );
  X_AND2   \BAR0/BR-15-8/$1I2989  (
    .I0(AD12),
    .I1(CFG13),
    .O(\BAR0/BR-15-8/IN4 )
  );
  X_AND2   \BAR0/BR-15-8/A2  (
    .I0(\BAR0/BR-15-8/EQ4 ),
    .I1(\BAR0/BR-15-8/EQ5 ),
    .O(\BAR0/BR-15-8/EQ54_5613 )
  );
  X_MUX2   \BAR0/BR-15-8/$1I2986  (
    .IB(\BAR0/BR-15-8/$1N2992 ),
    .IA(\BAR0/BR-15-8/$1N2910 ),
    .O(\BAR0/$1N3368 ),
    .SEL(\BAR0/BR-15-8/EQ76_5616 )
  );
  X_MUX2   \BAR0/BR-15-8/$1I2985  (
    .IB(\BAR0/BR-15-8/$1N2993 ),
    .IA(\BAR0/BR-15-8/$1N2911 ),
    .O(\BAR0/BR-15-8/$1N2992 ),
    .SEL(\BAR0/BR-15-8/EQ54_5613 )
  );
  X_AND2   \BAR0/BR-15-8/A3  (
    .I0(\BAR0/BR-15-8/EQ6 ),
    .I1(\BAR0/BR-15-8/EQ7 ),
    .O(\BAR0/BR-15-8/EQ76_5616 )
  );
  X_XOR2   \BAR0/BR-15-8/X4  (
    .I0(\BAR0/BR-15-8/IN4 ),
    .I1(\0BR12 ),
    .O(\NlwInverterSignal_BAR0/BR-15-8/X4/O )
  );
  X_XOR2   \BAR0/BR-15-8/X6  (
    .I0(\BAR0/BR-15-8/IN6 ),
    .I1(\0BR14 ),
    .O(\NlwInverterSignal_BAR0/BR-15-8/X6/O )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR0/BR-15-8/Q4  (
    .CE(CE4_1),
    .CLK(CLK),
    .I(AD12),
    .O(\BAR0/BR-15-8/RAWQ4 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR0/BR-15-8/Q5  (
    .CE(CE4_1),
    .CLK(CLK),
    .I(AD13),
    .O(\BAR0/BR-15-8/RAWQ5 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR0/BR-15-8/Q6  (
    .CE(CE4_1),
    .CLK(CLK),
    .I(AD14),
    .O(\BAR0/BR-15-8/RAWQ6 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR0/BR-15-8/Q7  (
    .CE(CE4_1),
    .CLK(CLK),
    .I(AD15),
    .O(\BAR0/BR-15-8/RAWQ7 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND2   \BAR0/BR-15-8/$1I2960  (
    .I0(AD15),
    .I1(CFG16),
    .O(\BAR0/BR-15-8/IN7 )
  );
  X_AND2   \BAR0/BR-15-8/$1I2959  (
    .I0(CFG16),
    .I1(\BAR0/BR-15-8/RAWQ7 ),
    .O(\0BR15 )
  );
  X_AND2   \BAR0/BR-15-8/$1I2958  (
    .I0(CFG13),
    .I1(\BAR0/BR-15-8/RAWQ4 ),
    .O(\0BR12 )
  );
  X_AND2   \BAR0/BR-15-8/$1I2957  (
    .I0(CFG14),
    .I1(\BAR0/BR-15-8/RAWQ5 ),
    .O(\0BR13 )
  );
  X_AND2   \BAR0/BR-15-8/$1I2956  (
    .I0(AD13),
    .I1(CFG14),
    .O(\BAR0/BR-15-8/IN5 )
  );
  X_AND2   \BAR0/BR-15-8/$1I2955  (
    .I0(AD14),
    .I1(CFG15),
    .O(\BAR0/BR-15-8/IN6 )
  );
  X_AND2   \BAR0/BR-15-8/$1I2954  (
    .I0(CFG15),
    .I1(\BAR0/BR-15-8/RAWQ6 ),
    .O(\0BR14 )
  );
  X_XOR2   \BAR0/BR-15-8/X7  (
    .I0(\BAR0/BR-15-8/IN7 ),
    .I1(\0BR15 ),
    .O(\NlwInverterSignal_BAR0/BR-15-8/X7/O )
  );
  X_XOR2   \BAR0/BR-15-8/X5  (
    .I0(\BAR0/BR-15-8/IN5 ),
    .I1(\0BR13 ),
    .O(\NlwInverterSignal_BAR0/BR-15-8/X5/O )
  );
  X_ZERO   \BAR0/BR-15-8/$1I2909/$1I2218  (
    .O(\BAR0/BR-15-8/$1I2909/$1N2216 )
  );
  X_BUF   \BAR0/BR-15-8/$1I2909/L  (
    .I(\BAR0/BR-15-8/$1I2909/$1N2216 ),
    .O(\BAR0/BR-15-8/$1N2910 )
  );
  X_ZERO   \BAR0/BR-15-8/$1I2990/$1I2218  (
    .O(\BAR0/BR-15-8/$1I2990/$1N2216 )
  );
  X_BUF   \BAR0/BR-15-8/$1I2990/L  (
    .I(\BAR0/BR-15-8/$1I2990/$1N2216 ),
    .O(\BAR0/BR-15-8/$1N2911 )
  );
  X_ZERO   \BAR0/BR-15-8/$1I3091/$1I2218  (
    .O(\BAR0/BR-15-8/$1I3091/$1N2216 )
  );
  X_BUF   \BAR0/BR-15-8/$1I3091/L  (
    .I(\BAR0/BR-15-8/$1I3091/$1N2216 ),
    .O(\BAR0/BR-15-8/$1N3110 )
  );
  X_ZERO   \BAR0/BR-15-8/$1I3096/$1I2218  (
    .O(\BAR0/BR-15-8/$1I3096/$1N2216 )
  );
  X_BUF   \BAR0/BR-15-8/$1I3096/L  (
    .I(\BAR0/BR-15-8/$1I3096/$1N2216 ),
    .O(\BAR0/BR-15-8/$1N3111 )
  );
  X_INV   \BAR0/BR-CMD/$1I228  (
    .I(EX),
    .O(\BAR0/BR-CMD/EX_N )
  );
  X_AND3   \BAR0/BR-CMD/$1I194  (
    .I0(\NlwInverterSignal_BAR0/BR-CMD/$1I194/I0 ),
    .I1(CBE_IN3),
    .I2(CBE_IN2),
    .O(\BAR0/BR-CMD/$1N195 )
  );
  X_OR2   \BAR0/BR-CMD/$1I193  (
    .I0(\BAR0/BR-CMD/$1N195 ),
    .I1(\BAR0/BR-CMD/$1N201 ),
    .O(\BAR0/BR-CMD/MEM_5666 )
  );
  X_AND2   \BAR0/BR-CMD/$1I192  (
    .I0(CBE_IN2),
    .I1(CBE_IN1),
    .O(\BAR0/BR-CMD/$1N201 )
  );
  X_AND3   \BAR0/BR-CMD/$1I173  (
    .I0(\NlwInverterSignal_BAR0/BR-CMD/$1I173/I0 ),
    .I1(\NlwInverterSignal_BAR0/BR-CMD/$1I173/I1 ),
    .I2(CBE_IN1),
    .O(\BAR0/BR-CMD/IO_5663 )
  );
  X_MUX2   \BAR0/BR-CMD/$1I157  (
    .IB(\BAR0/$1N3380 ),
    .IA(\BAR0/BR-CMD/$1N144 ),
    .O(\BAR0/MATCH ),
    .SEL(\BAR0/BR-CMD/SEL )
  );
  X_AND2   \BAR0/BR-CMD/$1I117  (
    .I0(\NlwInverterSignal_BAR0/BR-CMD/$1I117/I0 ),
    .I1(CFG35),
    .O(\0BR2 )
  );
  X_AND2   \BAR0/BR-CMD/$1I110  (
    .I0(\NlwInverterSignal_BAR0/BR-CMD/$1I110/I0 ),
    .I1(CFG34),
    .O(\0BR1 )
  );
  X_BUF   \BAR0/BR-CMD/$1I109  (
    .I(CFG36),
    .O(\0BR0 )
  );
  X_AND2   \BAR0/BR-CMD/$1I100  (
    .I0(\NlwInverterSignal_BAR0/BR-CMD/$1I100/I0 ),
    .I1(CFG33),
    .O(\0BR3 )
  );
  X_ZERO   \BAR0/BR-CMD/$1I143/$1I2218  (
    .O(\BAR0/BR-CMD/$1I143/$1N2216 )
  );
  X_BUF   \BAR0/BR-CMD/$1I143/L  (
    .I(\BAR0/BR-CMD/$1I143/$1N2216 ),
    .O(\BAR0/BR-CMD/$1N144 )
  );
  X_OR2   \BAR0/BR-CMD/$1I223/$1I38  (
    .I0(\BAR0/BR-CMD/$1I223/M1 ),
    .I1(\BAR0/BR-CMD/$1I223/M0 ),
    .O(\BAR0/BR-CMD/SEL )
  );
  X_AND3   \BAR0/BR-CMD/$1I223/$1I31  (
    .I0(\NlwInverterSignal_BAR0/BR-CMD/$1I223/$1I31/I0 ),
    .I1(\BAR0/BR-CMD/EX_N ),
    .I2(\BAR0/BR-CMD/MEM_5666 ),
    .O(\BAR0/BR-CMD/$1I223/M0 )
  );
  X_AND3   \BAR0/BR-CMD/$1I223/$1I30  (
    .I0(\BAR0/BR-CMD/IO_5663 ),
    .I1(\BAR0/BR-CMD/EX_N ),
    .I2(CFG36),
    .O(\BAR0/BR-CMD/$1I223/M1 )
  );
  X_MUX2   \BAR0/BR-7-4/$1I2695  (
    .IB(CFG0),
    .IA(\BAR0/BR-7-4/$1N2701 ),
    .O(\BAR0/BR-7-4/$1N2697 ),
    .SEL(\BAR0/BR-7-4/EQ54_5702 )
  );
  X_MUX2   \BAR0/BR-7-4/$1I2694  (
    .IB(\BAR0/BR-7-4/$1N2697 ),
    .IA(\BAR0/BR-7-4/$1N2706 ),
    .O(\BAR0/$1N3366 ),
    .SEL(\BAR0/BR-7-4/EQ76_5701 )
  );
  X_AND2   \BAR0/BR-7-4/$1I2676  (
    .I0(AD4),
    .I1(CFG5),
    .O(\BAR0/BR-7-4/IN4 )
  );
  X_AND2   \BAR0/BR-7-4/$1I2672  (
    .I0(AD5),
    .I1(CFG6),
    .O(\BAR0/BR-7-4/IN5 )
  );
  X_AND2   \BAR0/BR-7-4/$1I2668  (
    .I0(AD6),
    .I1(CFG7),
    .O(\BAR0/BR-7-4/IN6 )
  );
  X_AND2   \BAR0/BR-7-4/$1I2664  (
    .I0(AD7),
    .I1(CFG8),
    .O(\BAR0/BR-7-4/IN7 )
  );
  X_AND2   \BAR0/BR-7-4/$1I2616  (
    .I0(CFG5),
    .I1(\BAR0/BR-7-4/RAWQ4 ),
    .O(\0BR4 )
  );
  X_AND2   \BAR0/BR-7-4/$1I2612  (
    .I0(CFG6),
    .I1(\BAR0/BR-7-4/RAWQ5 ),
    .O(\0BR5 )
  );
  X_AND2   \BAR0/BR-7-4/$1I2608  (
    .I0(CFG7),
    .I1(\BAR0/BR-7-4/RAWQ6 ),
    .O(\0BR6 )
  );
  X_AND2   \BAR0/BR-7-4/$1I2602  (
    .I0(CFG8),
    .I1(\BAR0/BR-7-4/RAWQ7 ),
    .O(\0BR7 )
  );
  X_AND2   \BAR0/BR-7-4/A2  (
    .I0(\BAR0/BR-7-4/EQ4 ),
    .I1(\BAR0/BR-7-4/EQ5 ),
    .O(\BAR0/BR-7-4/EQ54_5702 )
  );
  X_AND2   \BAR0/BR-7-4/A3  (
    .I0(\BAR0/BR-7-4/EQ6 ),
    .I1(\BAR0/BR-7-4/EQ7 ),
    .O(\BAR0/BR-7-4/EQ76_5701 )
  );
  X_XOR2   \BAR0/BR-7-4/X7  (
    .I0(\BAR0/BR-7-4/IN7 ),
    .I1(\0BR7 ),
    .O(\NlwInverterSignal_BAR0/BR-7-4/X7/O )
  );
  X_XOR2   \BAR0/BR-7-4/X6  (
    .I0(\BAR0/BR-7-4/IN6 ),
    .I1(\0BR6 ),
    .O(\NlwInverterSignal_BAR0/BR-7-4/X6/O )
  );
  X_XOR2   \BAR0/BR-7-4/X5  (
    .I0(\BAR0/BR-7-4/IN5 ),
    .I1(\0BR5 ),
    .O(\NlwInverterSignal_BAR0/BR-7-4/X5/O )
  );
  X_XOR2   \BAR0/BR-7-4/X4  (
    .I0(\BAR0/BR-7-4/IN4 ),
    .I1(\0BR4 ),
    .O(\NlwInverterSignal_BAR0/BR-7-4/X4/O )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR0/BR-7-4/Q7  (
    .CE(CE4_0),
    .CLK(CLK),
    .I(AD7),
    .O(\BAR0/BR-7-4/RAWQ7 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR0/BR-7-4/Q6  (
    .CE(CE4_0),
    .CLK(CLK),
    .I(AD6),
    .O(\BAR0/BR-7-4/RAWQ6 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR0/BR-7-4/Q5  (
    .CE(CE4_0),
    .CLK(CLK),
    .I(AD5),
    .O(\BAR0/BR-7-4/RAWQ5 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR0/BR-7-4/Q4  (
    .CE(CE4_0),
    .CLK(CLK),
    .I(AD4),
    .O(\BAR0/BR-7-4/RAWQ4 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_ZERO   \BAR0/BR-7-4/$1I2700/$1I2218  (
    .O(\BAR0/BR-7-4/$1I2700/$1N2216 )
  );
  X_BUF   \BAR0/BR-7-4/$1I2700/L  (
    .I(\BAR0/BR-7-4/$1I2700/$1N2216 ),
    .O(\BAR0/BR-7-4/$1N2701 )
  );
  X_ZERO   \BAR0/BR-7-4/$1I2705/$1I2218  (
    .O(\BAR0/BR-7-4/$1I2705/$1N2216 )
  );
  X_BUF   \BAR0/BR-7-4/$1I2705/L  (
    .I(\BAR0/BR-7-4/$1I2705/$1N2216 ),
    .O(\BAR0/BR-7-4/$1N2706 )
  );
  X_OR2   \BAR0/$1I3440/$1I38  (
    .I0(\BAR0/$1I3440/M1 ),
    .I1(\BAR0/$1I3440/M0 ),
    .O(\BAR0/CSREN32 )
  );
  X_AND3   \BAR0/$1I3440/$1I31  (
    .I0(\NlwInverterSignal_BAR0/$1I3440/$1I31/I0 ),
    .I1(CFG0),
    .I2(NlwRenamedSig_OI_CSR1),
    .O(\BAR0/$1I3440/M0 )
  );
  X_AND3   \BAR0/$1I3440/$1I30  (
    .I0(NlwRenamedSig_OI_CSR0),
    .I1(CFG0),
    .I2(CFG36),
    .O(\BAR0/$1I3440/M1 )
  );
  X_OR2   \BAR0/$1I3453/$1I38  (
    .I0(\BAR0/$1I3453/M1 ),
    .I1(\BAR0/$1I3453/M0 ),
    .O(\BAR0/CSREN64 )
  );
  X_AND3   \BAR0/$1I3453/$1I31  (
    .I0(\NlwInverterSignal_BAR0/$1I3453/$1I31/I0 ),
    .I1(CFG0),
    .I2(NlwRenamedSig_OI_CSR1),
    .O(\BAR0/$1I3453/M0 )
  );
  X_AND3   \BAR0/$1I3453/$1I30  (
    .I0(\BAR0/$1N3458 ),
    .I1(CFG0),
    .I2(CFG36),
    .O(\BAR0/$1I3453/M1 )
  );
  X_ZERO   \BAR0/$1I3468/$1I2218  (
    .O(\BAR0/$1I3468/$1N2216 )
  );
  X_BUF   \BAR0/$1I3468/L  (
    .I(\BAR0/$1I3468/$1N2216 ),
    .O(\BAR0/$1N3458 )
  );
  X_ONE   \BAR0/$1I3469/$1I2220  (
    .O(\BAR0/$1I3469/$1N2216 )
  );
  X_BUF   \BAR0/$1I3469/H  (
    .I(\BAR0/$1I3469/$1N2216 ),
    .O(\BAR0/ENABLE32 )
  );
  X_ONE   \BAR0/$2I3304/$1I2220  (
    .O(\BAR0/$2I3304/$1N2216 )
  );
  X_BUF   \BAR0/$2I3304/H  (
    .I(\BAR0/$2I3304/$1N2216 ),
    .O(\BAR0/ENABLENL )
  );
  X_OR2   \BAR0/$2I3321/$1I38  (
    .I0(\BAR0/$2I3321/M1 ),
    .I1(\BAR0/$2I3321/M0 ),
    .O(\BAR0/CSRENNL )
  );
  X_AND3   \BAR0/$2I3321/$1I31  (
    .I0(\NlwInverterSignal_BAR0/$2I3321/$1I31/I0 ),
    .I1(CFG0),
    .I2(NlwRenamedSig_OI_CSR1),
    .O(\BAR0/$2I3321/M0 )
  );
  X_AND3   \BAR0/$2I3321/$1I30  (
    .I0(NlwRenamedSig_OI_CSR0),
    .I1(CFG0),
    .I2(CFG36),
    .O(\BAR0/$2I3321/M1 )
  );
  X_AND4   \BAR1/$2I3324  (
    .I0(\BAR1/CSRENNL ),
    .I1(\BAR1/MATCH ),
    .I2(ADDR_VLD1),
    .I3(\BAR1/ENABLENL ),
    .O(\BAR1/NS_HITNL )
  );
  X_INV   \BAR1/$2I3284  (
    .I(CFG73),
    .O(\BAR1/NL_CE )
  );
  X_AND2   \BAR1/$2I3275  (
    .I0(\TSTOP_I- ),
    .I1(\BAR1/$2N3280 ),
    .O(\BAR1/NS_NL_MEM )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR1/NL  (
    .CE(\BAR1/NL_CE ),
    .CLK(CLK),
    .I(\BAR1/NS_NL_MEM ),
    .O(NL_MEM1),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_OR2   \BAR1/$2I3268  (
    .I0(\BAR1/$2N3273 ),
    .I1(NL_MEM1),
    .O(\BAR1/$2N3280 )
  );
  X_AND2   \BAR1/$2I3267  (
    .I0(\BAR1/UNALIGN ),
    .I1(\BAR1/NS_HITNL ),
    .O(\BAR1/$2N3273 )
  );
  X_OR2   \BAR1/$2I3263  (
    .I0(AD1),
    .I1(AD0),
    .O(\BAR1/UNALIGN )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR1/EQ64  (
    .CE(VCC),
    .CLK(CLK),
    .I(NS_BH64_1),
    .O(BH64_1),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR1/EQ32  (
    .CE(VCC),
    .CLK(CLK),
    .I(NS_BASE_HIT1),
    .O(NlwRenamedSig_OI_BASE_HIT1),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND4   \BAR1/$1I3455  (
    .I0(\BAR1/CSREN64 ),
    .I1(\BAR1/MATCH ),
    .I2(ADDR_VLD64),
    .I3(CFG242),
    .O(NS_BH64_1)
  );
  X_AND4   \BAR1/$1I3437  (
    .I0(\BAR1/CSREN32 ),
    .I1(\BAR1/MATCH ),
    .I2(ADDR_VLD1),
    .I3(\BAR1/ENABLE32 ),
    .O(NS_BASE_HIT1)
  );
  X_MUX2   \BAR1/BR-31-24/$1I3094  (
    .IB(\BAR1/$1N3369 ),
    .IA(\BAR1/BR-31-24/$1N3110 ),
    .O(\BAR1/BR-31-24/$1N3099 ),
    .SEL(\BAR1/BR-31-24/EQ10_5938 )
  );
  X_MUX2   \BAR1/BR-31-24/$1I3093  (
    .IB(\BAR1/BR-31-24/$1N3099 ),
    .IA(\BAR1/BR-31-24/$1N3111 ),
    .O(\BAR1/BR-31-24/$1N2993 ),
    .SEL(\BAR1/BR-31-24/EQ32_5941 )
  );
  X_XOR2   \BAR1/BR-31-24/X1  (
    .I0(\BAR1/BR-31-24/IN1 ),
    .I1(\1BR25 ),
    .O(\NlwInverterSignal_BAR1/BR-31-24/X1/O )
  );
  X_XOR2   \BAR1/BR-31-24/X3  (
    .I0(\BAR1/BR-31-24/IN3 ),
    .I1(\1BR27 ),
    .O(\NlwInverterSignal_BAR1/BR-31-24/X3/O )
  );
  X_AND2   \BAR1/BR-31-24/$1I3014  (
    .I0(CFG64),
    .I1(\BAR1/BR-31-24/RAWQ2 ),
    .O(\1BR26 )
  );
  X_AND2   \BAR1/BR-31-24/$1I3013  (
    .I0(AD26),
    .I1(CFG64),
    .O(\BAR1/BR-31-24/IN2 )
  );
  X_AND2   \BAR1/BR-31-24/$1I3012  (
    .I0(AD25),
    .I1(CFG63),
    .O(\BAR1/BR-31-24/IN1 )
  );
  X_AND2   \BAR1/BR-31-24/$1I3011  (
    .I0(CFG63),
    .I1(\BAR1/BR-31-24/RAWQ1 ),
    .O(\1BR25 )
  );
  X_AND2   \BAR1/BR-31-24/$1I3010  (
    .I0(CFG62),
    .I1(\BAR1/BR-31-24/RAWQ0 ),
    .O(\1BR24 )
  );
  X_AND2   \BAR1/BR-31-24/$1I3009  (
    .I0(CFG65),
    .I1(\BAR1/BR-31-24/RAWQ3 ),
    .O(\1BR27 )
  );
  X_AND2   \BAR1/BR-31-24/$1I3008  (
    .I0(AD27),
    .I1(CFG65),
    .O(\BAR1/BR-31-24/IN3 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR1/BR-31-24/Q3  (
    .CE(CE5_3),
    .CLK(CLK),
    .I(AD27),
    .O(\BAR1/BR-31-24/RAWQ3 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR1/BR-31-24/Q2  (
    .CE(CE5_3),
    .CLK(CLK),
    .I(AD26),
    .O(\BAR1/BR-31-24/RAWQ2 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR1/BR-31-24/Q1  (
    .CE(CE5_3),
    .CLK(CLK),
    .I(AD25),
    .O(\BAR1/BR-31-24/RAWQ1 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR1/BR-31-24/Q0  (
    .CE(CE5_3),
    .CLK(CLK),
    .I(AD24),
    .O(\BAR1/BR-31-24/RAWQ0 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \BAR1/BR-31-24/X2  (
    .I0(\BAR1/BR-31-24/IN2 ),
    .I1(\1BR26 ),
    .O(\NlwInverterSignal_BAR1/BR-31-24/X2/O )
  );
  X_XOR2   \BAR1/BR-31-24/X0  (
    .I0(\BAR1/BR-31-24/IN0 ),
    .I1(\1BR24 ),
    .O(\NlwInverterSignal_BAR1/BR-31-24/X0/O )
  );
  X_AND2   \BAR1/BR-31-24/A1  (
    .I0(\BAR1/BR-31-24/EQ2 ),
    .I1(\BAR1/BR-31-24/EQ3 ),
    .O(\BAR1/BR-31-24/EQ32_5941 )
  );
  X_AND2   \BAR1/BR-31-24/A0  (
    .I0(\BAR1/BR-31-24/EQ0 ),
    .I1(\BAR1/BR-31-24/EQ1 ),
    .O(\BAR1/BR-31-24/EQ10_5938 )
  );
  X_AND2   \BAR1/BR-31-24/$1I2999  (
    .I0(AD24),
    .I1(CFG62),
    .O(\BAR1/BR-31-24/IN0 )
  );
  X_AND2   \BAR1/BR-31-24/$1I2989  (
    .I0(AD28),
    .I1(CFG66),
    .O(\BAR1/BR-31-24/IN4 )
  );
  X_AND2   \BAR1/BR-31-24/A2  (
    .I0(\BAR1/BR-31-24/EQ4 ),
    .I1(\BAR1/BR-31-24/EQ5 ),
    .O(\BAR1/BR-31-24/EQ54_5928 )
  );
  X_MUX2   \BAR1/BR-31-24/$1I2986  (
    .IB(\BAR1/BR-31-24/$1N2992 ),
    .IA(\BAR1/BR-31-24/$1N2910 ),
    .O(\BAR1/$1N3380 ),
    .SEL(\BAR1/BR-31-24/EQ76_5931 )
  );
  X_MUX2   \BAR1/BR-31-24/$1I2985  (
    .IB(\BAR1/BR-31-24/$1N2993 ),
    .IA(\BAR1/BR-31-24/$1N2911 ),
    .O(\BAR1/BR-31-24/$1N2992 ),
    .SEL(\BAR1/BR-31-24/EQ54_5928 )
  );
  X_AND2   \BAR1/BR-31-24/A3  (
    .I0(\BAR1/BR-31-24/EQ6 ),
    .I1(\BAR1/BR-31-24/EQ7 ),
    .O(\BAR1/BR-31-24/EQ76_5931 )
  );
  X_XOR2   \BAR1/BR-31-24/X4  (
    .I0(\BAR1/BR-31-24/IN4 ),
    .I1(\1BR28 ),
    .O(\NlwInverterSignal_BAR1/BR-31-24/X4/O )
  );
  X_XOR2   \BAR1/BR-31-24/X6  (
    .I0(\BAR1/BR-31-24/IN6 ),
    .I1(\1BR30 ),
    .O(\NlwInverterSignal_BAR1/BR-31-24/X6/O )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR1/BR-31-24/Q4  (
    .CE(CE5_3),
    .CLK(CLK),
    .I(AD28),
    .O(\BAR1/BR-31-24/RAWQ4 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR1/BR-31-24/Q5  (
    .CE(CE5_3),
    .CLK(CLK),
    .I(AD29),
    .O(\BAR1/BR-31-24/RAWQ5 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR1/BR-31-24/Q6  (
    .CE(CE5_3),
    .CLK(CLK),
    .I(AD30),
    .O(\BAR1/BR-31-24/RAWQ6 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR1/BR-31-24/Q7  (
    .CE(CE5_3),
    .CLK(CLK),
    .I(AD31),
    .O(\BAR1/BR-31-24/RAWQ7 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND2   \BAR1/BR-31-24/$1I2960  (
    .I0(AD31),
    .I1(CFG69),
    .O(\BAR1/BR-31-24/IN7 )
  );
  X_AND2   \BAR1/BR-31-24/$1I2959  (
    .I0(CFG69),
    .I1(\BAR1/BR-31-24/RAWQ7 ),
    .O(\1BR31 )
  );
  X_AND2   \BAR1/BR-31-24/$1I2958  (
    .I0(CFG66),
    .I1(\BAR1/BR-31-24/RAWQ4 ),
    .O(\1BR28 )
  );
  X_AND2   \BAR1/BR-31-24/$1I2957  (
    .I0(CFG67),
    .I1(\BAR1/BR-31-24/RAWQ5 ),
    .O(\1BR29 )
  );
  X_AND2   \BAR1/BR-31-24/$1I2956  (
    .I0(AD29),
    .I1(CFG67),
    .O(\BAR1/BR-31-24/IN5 )
  );
  X_AND2   \BAR1/BR-31-24/$1I2955  (
    .I0(AD30),
    .I1(CFG68),
    .O(\BAR1/BR-31-24/IN6 )
  );
  X_AND2   \BAR1/BR-31-24/$1I2954  (
    .I0(CFG68),
    .I1(\BAR1/BR-31-24/RAWQ6 ),
    .O(\1BR30 )
  );
  X_XOR2   \BAR1/BR-31-24/X7  (
    .I0(\BAR1/BR-31-24/IN7 ),
    .I1(\1BR31 ),
    .O(\NlwInverterSignal_BAR1/BR-31-24/X7/O )
  );
  X_XOR2   \BAR1/BR-31-24/X5  (
    .I0(\BAR1/BR-31-24/IN5 ),
    .I1(\1BR29 ),
    .O(\NlwInverterSignal_BAR1/BR-31-24/X5/O )
  );
  X_ZERO   \BAR1/BR-31-24/$1I2909/$1I2218  (
    .O(\BAR1/BR-31-24/$1I2909/$1N2216 )
  );
  X_BUF   \BAR1/BR-31-24/$1I2909/L  (
    .I(\BAR1/BR-31-24/$1I2909/$1N2216 ),
    .O(\BAR1/BR-31-24/$1N2910 )
  );
  X_ZERO   \BAR1/BR-31-24/$1I2990/$1I2218  (
    .O(\BAR1/BR-31-24/$1I2990/$1N2216 )
  );
  X_BUF   \BAR1/BR-31-24/$1I2990/L  (
    .I(\BAR1/BR-31-24/$1I2990/$1N2216 ),
    .O(\BAR1/BR-31-24/$1N2911 )
  );
  X_ZERO   \BAR1/BR-31-24/$1I3091/$1I2218  (
    .O(\BAR1/BR-31-24/$1I3091/$1N2216 )
  );
  X_BUF   \BAR1/BR-31-24/$1I3091/L  (
    .I(\BAR1/BR-31-24/$1I3091/$1N2216 ),
    .O(\BAR1/BR-31-24/$1N3110 )
  );
  X_ZERO   \BAR1/BR-31-24/$1I3096/$1I2218  (
    .O(\BAR1/BR-31-24/$1I3096/$1N2216 )
  );
  X_BUF   \BAR1/BR-31-24/$1I3096/L  (
    .I(\BAR1/BR-31-24/$1I3096/$1N2216 ),
    .O(\BAR1/BR-31-24/$1N3111 )
  );
  X_MUX2   \BAR1/BR-23-16/$1I3094  (
    .IB(\BAR1/$1N3368 ),
    .IA(\BAR1/BR-23-16/$1N3110 ),
    .O(\BAR1/BR-23-16/$1N3099 ),
    .SEL(\BAR1/BR-23-16/EQ10_6010 )
  );
  X_MUX2   \BAR1/BR-23-16/$1I3093  (
    .IB(\BAR1/BR-23-16/$1N3099 ),
    .IA(\BAR1/BR-23-16/$1N3111 ),
    .O(\BAR1/BR-23-16/$1N2993 ),
    .SEL(\BAR1/BR-23-16/EQ32_6013 )
  );
  X_XOR2   \BAR1/BR-23-16/X1  (
    .I0(\BAR1/BR-23-16/IN1 ),
    .I1(\1BR17 ),
    .O(\NlwInverterSignal_BAR1/BR-23-16/X1/O )
  );
  X_XOR2   \BAR1/BR-23-16/X3  (
    .I0(\BAR1/BR-23-16/IN3 ),
    .I1(\1BR19 ),
    .O(\NlwInverterSignal_BAR1/BR-23-16/X3/O )
  );
  X_AND2   \BAR1/BR-23-16/$1I3014  (
    .I0(CFG56),
    .I1(\BAR1/BR-23-16/RAWQ2 ),
    .O(\1BR18 )
  );
  X_AND2   \BAR1/BR-23-16/$1I3013  (
    .I0(AD18),
    .I1(CFG56),
    .O(\BAR1/BR-23-16/IN2 )
  );
  X_AND2   \BAR1/BR-23-16/$1I3012  (
    .I0(AD17),
    .I1(CFG55),
    .O(\BAR1/BR-23-16/IN1 )
  );
  X_AND2   \BAR1/BR-23-16/$1I3011  (
    .I0(CFG55),
    .I1(\BAR1/BR-23-16/RAWQ1 ),
    .O(\1BR17 )
  );
  X_AND2   \BAR1/BR-23-16/$1I3010  (
    .I0(CFG54),
    .I1(\BAR1/BR-23-16/RAWQ0 ),
    .O(\1BR16 )
  );
  X_AND2   \BAR1/BR-23-16/$1I3009  (
    .I0(CFG57),
    .I1(\BAR1/BR-23-16/RAWQ3 ),
    .O(\1BR19 )
  );
  X_AND2   \BAR1/BR-23-16/$1I3008  (
    .I0(AD19),
    .I1(CFG57),
    .O(\BAR1/BR-23-16/IN3 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR1/BR-23-16/Q3  (
    .CE(CE5_2),
    .CLK(CLK),
    .I(AD19),
    .O(\BAR1/BR-23-16/RAWQ3 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR1/BR-23-16/Q2  (
    .CE(CE5_2),
    .CLK(CLK),
    .I(AD18),
    .O(\BAR1/BR-23-16/RAWQ2 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR1/BR-23-16/Q1  (
    .CE(CE5_2),
    .CLK(CLK),
    .I(AD17),
    .O(\BAR1/BR-23-16/RAWQ1 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR1/BR-23-16/Q0  (
    .CE(CE5_2),
    .CLK(CLK),
    .I(AD16),
    .O(\BAR1/BR-23-16/RAWQ0 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \BAR1/BR-23-16/X2  (
    .I0(\BAR1/BR-23-16/IN2 ),
    .I1(\1BR18 ),
    .O(\NlwInverterSignal_BAR1/BR-23-16/X2/O )
  );
  X_XOR2   \BAR1/BR-23-16/X0  (
    .I0(\BAR1/BR-23-16/IN0 ),
    .I1(\1BR16 ),
    .O(\NlwInverterSignal_BAR1/BR-23-16/X0/O )
  );
  X_AND2   \BAR1/BR-23-16/A1  (
    .I0(\BAR1/BR-23-16/EQ2 ),
    .I1(\BAR1/BR-23-16/EQ3 ),
    .O(\BAR1/BR-23-16/EQ32_6013 )
  );
  X_AND2   \BAR1/BR-23-16/A0  (
    .I0(\BAR1/BR-23-16/EQ0 ),
    .I1(\BAR1/BR-23-16/EQ1 ),
    .O(\BAR1/BR-23-16/EQ10_6010 )
  );
  X_AND2   \BAR1/BR-23-16/$1I2999  (
    .I0(AD16),
    .I1(CFG54),
    .O(\BAR1/BR-23-16/IN0 )
  );
  X_AND2   \BAR1/BR-23-16/$1I2989  (
    .I0(AD20),
    .I1(CFG58),
    .O(\BAR1/BR-23-16/IN4 )
  );
  X_AND2   \BAR1/BR-23-16/A2  (
    .I0(\BAR1/BR-23-16/EQ4 ),
    .I1(\BAR1/BR-23-16/EQ5 ),
    .O(\BAR1/BR-23-16/EQ54_6000 )
  );
  X_MUX2   \BAR1/BR-23-16/$1I2986  (
    .IB(\BAR1/BR-23-16/$1N2992 ),
    .IA(\BAR1/BR-23-16/$1N2910 ),
    .O(\BAR1/$1N3369 ),
    .SEL(\BAR1/BR-23-16/EQ76_6003 )
  );
  X_MUX2   \BAR1/BR-23-16/$1I2985  (
    .IB(\BAR1/BR-23-16/$1N2993 ),
    .IA(\BAR1/BR-23-16/$1N2911 ),
    .O(\BAR1/BR-23-16/$1N2992 ),
    .SEL(\BAR1/BR-23-16/EQ54_6000 )
  );
  X_AND2   \BAR1/BR-23-16/A3  (
    .I0(\BAR1/BR-23-16/EQ6 ),
    .I1(\BAR1/BR-23-16/EQ7 ),
    .O(\BAR1/BR-23-16/EQ76_6003 )
  );
  X_XOR2   \BAR1/BR-23-16/X4  (
    .I0(\BAR1/BR-23-16/IN4 ),
    .I1(\1BR20 ),
    .O(\NlwInverterSignal_BAR1/BR-23-16/X4/O )
  );
  X_XOR2   \BAR1/BR-23-16/X6  (
    .I0(\BAR1/BR-23-16/IN6 ),
    .I1(\1BR22 ),
    .O(\NlwInverterSignal_BAR1/BR-23-16/X6/O )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR1/BR-23-16/Q4  (
    .CE(CE5_2),
    .CLK(CLK),
    .I(AD20),
    .O(\BAR1/BR-23-16/RAWQ4 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR1/BR-23-16/Q5  (
    .CE(CE5_2),
    .CLK(CLK),
    .I(AD21),
    .O(\BAR1/BR-23-16/RAWQ5 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR1/BR-23-16/Q6  (
    .CE(CE5_2),
    .CLK(CLK),
    .I(AD22),
    .O(\BAR1/BR-23-16/RAWQ6 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR1/BR-23-16/Q7  (
    .CE(CE5_2),
    .CLK(CLK),
    .I(AD23),
    .O(\BAR1/BR-23-16/RAWQ7 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND2   \BAR1/BR-23-16/$1I2960  (
    .I0(AD23),
    .I1(CFG61),
    .O(\BAR1/BR-23-16/IN7 )
  );
  X_AND2   \BAR1/BR-23-16/$1I2959  (
    .I0(CFG61),
    .I1(\BAR1/BR-23-16/RAWQ7 ),
    .O(\1BR23 )
  );
  X_AND2   \BAR1/BR-23-16/$1I2958  (
    .I0(CFG58),
    .I1(\BAR1/BR-23-16/RAWQ4 ),
    .O(\1BR20 )
  );
  X_AND2   \BAR1/BR-23-16/$1I2957  (
    .I0(CFG59),
    .I1(\BAR1/BR-23-16/RAWQ5 ),
    .O(\1BR21 )
  );
  X_AND2   \BAR1/BR-23-16/$1I2956  (
    .I0(AD21),
    .I1(CFG59),
    .O(\BAR1/BR-23-16/IN5 )
  );
  X_AND2   \BAR1/BR-23-16/$1I2955  (
    .I0(AD22),
    .I1(CFG60),
    .O(\BAR1/BR-23-16/IN6 )
  );
  X_AND2   \BAR1/BR-23-16/$1I2954  (
    .I0(CFG60),
    .I1(\BAR1/BR-23-16/RAWQ6 ),
    .O(\1BR22 )
  );
  X_XOR2   \BAR1/BR-23-16/X7  (
    .I0(\BAR1/BR-23-16/IN7 ),
    .I1(\1BR23 ),
    .O(\NlwInverterSignal_BAR1/BR-23-16/X7/O )
  );
  X_XOR2   \BAR1/BR-23-16/X5  (
    .I0(\BAR1/BR-23-16/IN5 ),
    .I1(\1BR21 ),
    .O(\NlwInverterSignal_BAR1/BR-23-16/X5/O )
  );
  X_ZERO   \BAR1/BR-23-16/$1I2909/$1I2218  (
    .O(\BAR1/BR-23-16/$1I2909/$1N2216 )
  );
  X_BUF   \BAR1/BR-23-16/$1I2909/L  (
    .I(\BAR1/BR-23-16/$1I2909/$1N2216 ),
    .O(\BAR1/BR-23-16/$1N2910 )
  );
  X_ZERO   \BAR1/BR-23-16/$1I2990/$1I2218  (
    .O(\BAR1/BR-23-16/$1I2990/$1N2216 )
  );
  X_BUF   \BAR1/BR-23-16/$1I2990/L  (
    .I(\BAR1/BR-23-16/$1I2990/$1N2216 ),
    .O(\BAR1/BR-23-16/$1N2911 )
  );
  X_ZERO   \BAR1/BR-23-16/$1I3091/$1I2218  (
    .O(\BAR1/BR-23-16/$1I3091/$1N2216 )
  );
  X_BUF   \BAR1/BR-23-16/$1I3091/L  (
    .I(\BAR1/BR-23-16/$1I3091/$1N2216 ),
    .O(\BAR1/BR-23-16/$1N3110 )
  );
  X_ZERO   \BAR1/BR-23-16/$1I3096/$1I2218  (
    .O(\BAR1/BR-23-16/$1I3096/$1N2216 )
  );
  X_BUF   \BAR1/BR-23-16/$1I3096/L  (
    .I(\BAR1/BR-23-16/$1I3096/$1N2216 ),
    .O(\BAR1/BR-23-16/$1N3111 )
  );
  X_MUX2   \BAR1/BR-15-8/$1I3094  (
    .IB(\BAR1/$1N3366 ),
    .IA(\BAR1/BR-15-8/$1N3110 ),
    .O(\BAR1/BR-15-8/$1N3099 ),
    .SEL(\BAR1/BR-15-8/EQ10_6082 )
  );
  X_MUX2   \BAR1/BR-15-8/$1I3093  (
    .IB(\BAR1/BR-15-8/$1N3099 ),
    .IA(\BAR1/BR-15-8/$1N3111 ),
    .O(\BAR1/BR-15-8/$1N2993 ),
    .SEL(\BAR1/BR-15-8/EQ32_6085 )
  );
  X_XOR2   \BAR1/BR-15-8/X1  (
    .I0(\BAR1/BR-15-8/IN1 ),
    .I1(\1BR9 ),
    .O(\NlwInverterSignal_BAR1/BR-15-8/X1/O )
  );
  X_XOR2   \BAR1/BR-15-8/X3  (
    .I0(\BAR1/BR-15-8/IN3 ),
    .I1(\1BR11 ),
    .O(\NlwInverterSignal_BAR1/BR-15-8/X3/O )
  );
  X_AND2   \BAR1/BR-15-8/$1I3014  (
    .I0(CFG48),
    .I1(\BAR1/BR-15-8/RAWQ2 ),
    .O(\1BR10 )
  );
  X_AND2   \BAR1/BR-15-8/$1I3013  (
    .I0(AD10),
    .I1(CFG48),
    .O(\BAR1/BR-15-8/IN2 )
  );
  X_AND2   \BAR1/BR-15-8/$1I3012  (
    .I0(AD9),
    .I1(CFG47),
    .O(\BAR1/BR-15-8/IN1 )
  );
  X_AND2   \BAR1/BR-15-8/$1I3011  (
    .I0(CFG47),
    .I1(\BAR1/BR-15-8/RAWQ1 ),
    .O(\1BR9 )
  );
  X_AND2   \BAR1/BR-15-8/$1I3010  (
    .I0(CFG46),
    .I1(\BAR1/BR-15-8/RAWQ0 ),
    .O(\1BR8 )
  );
  X_AND2   \BAR1/BR-15-8/$1I3009  (
    .I0(CFG49),
    .I1(\BAR1/BR-15-8/RAWQ3 ),
    .O(\1BR11 )
  );
  X_AND2   \BAR1/BR-15-8/$1I3008  (
    .I0(AD11),
    .I1(CFG49),
    .O(\BAR1/BR-15-8/IN3 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR1/BR-15-8/Q3  (
    .CE(CE5_1),
    .CLK(CLK),
    .I(AD11),
    .O(\BAR1/BR-15-8/RAWQ3 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR1/BR-15-8/Q2  (
    .CE(CE5_1),
    .CLK(CLK),
    .I(AD10),
    .O(\BAR1/BR-15-8/RAWQ2 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR1/BR-15-8/Q1  (
    .CE(CE5_1),
    .CLK(CLK),
    .I(AD9),
    .O(\BAR1/BR-15-8/RAWQ1 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR1/BR-15-8/Q0  (
    .CE(CE5_1),
    .CLK(CLK),
    .I(AD8),
    .O(\BAR1/BR-15-8/RAWQ0 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \BAR1/BR-15-8/X2  (
    .I0(\BAR1/BR-15-8/IN2 ),
    .I1(\1BR10 ),
    .O(\NlwInverterSignal_BAR1/BR-15-8/X2/O )
  );
  X_XOR2   \BAR1/BR-15-8/X0  (
    .I0(\BAR1/BR-15-8/IN0 ),
    .I1(\1BR8 ),
    .O(\NlwInverterSignal_BAR1/BR-15-8/X0/O )
  );
  X_AND2   \BAR1/BR-15-8/A1  (
    .I0(\BAR1/BR-15-8/EQ2 ),
    .I1(\BAR1/BR-15-8/EQ3 ),
    .O(\BAR1/BR-15-8/EQ32_6085 )
  );
  X_AND2   \BAR1/BR-15-8/A0  (
    .I0(\BAR1/BR-15-8/EQ0 ),
    .I1(\BAR1/BR-15-8/EQ1 ),
    .O(\BAR1/BR-15-8/EQ10_6082 )
  );
  X_AND2   \BAR1/BR-15-8/$1I2999  (
    .I0(AD8),
    .I1(CFG46),
    .O(\BAR1/BR-15-8/IN0 )
  );
  X_AND2   \BAR1/BR-15-8/$1I2989  (
    .I0(AD12),
    .I1(CFG50),
    .O(\BAR1/BR-15-8/IN4 )
  );
  X_AND2   \BAR1/BR-15-8/A2  (
    .I0(\BAR1/BR-15-8/EQ4 ),
    .I1(\BAR1/BR-15-8/EQ5 ),
    .O(\BAR1/BR-15-8/EQ54_6072 )
  );
  X_MUX2   \BAR1/BR-15-8/$1I2986  (
    .IB(\BAR1/BR-15-8/$1N2992 ),
    .IA(\BAR1/BR-15-8/$1N2910 ),
    .O(\BAR1/$1N3368 ),
    .SEL(\BAR1/BR-15-8/EQ76_6075 )
  );
  X_MUX2   \BAR1/BR-15-8/$1I2985  (
    .IB(\BAR1/BR-15-8/$1N2993 ),
    .IA(\BAR1/BR-15-8/$1N2911 ),
    .O(\BAR1/BR-15-8/$1N2992 ),
    .SEL(\BAR1/BR-15-8/EQ54_6072 )
  );
  X_AND2   \BAR1/BR-15-8/A3  (
    .I0(\BAR1/BR-15-8/EQ6 ),
    .I1(\BAR1/BR-15-8/EQ7 ),
    .O(\BAR1/BR-15-8/EQ76_6075 )
  );
  X_XOR2   \BAR1/BR-15-8/X4  (
    .I0(\BAR1/BR-15-8/IN4 ),
    .I1(\1BR12 ),
    .O(\NlwInverterSignal_BAR1/BR-15-8/X4/O )
  );
  X_XOR2   \BAR1/BR-15-8/X6  (
    .I0(\BAR1/BR-15-8/IN6 ),
    .I1(\1BR14 ),
    .O(\NlwInverterSignal_BAR1/BR-15-8/X6/O )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR1/BR-15-8/Q4  (
    .CE(CE5_1),
    .CLK(CLK),
    .I(AD12),
    .O(\BAR1/BR-15-8/RAWQ4 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR1/BR-15-8/Q5  (
    .CE(CE5_1),
    .CLK(CLK),
    .I(AD13),
    .O(\BAR1/BR-15-8/RAWQ5 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR1/BR-15-8/Q6  (
    .CE(CE5_1),
    .CLK(CLK),
    .I(AD14),
    .O(\BAR1/BR-15-8/RAWQ6 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR1/BR-15-8/Q7  (
    .CE(CE5_1),
    .CLK(CLK),
    .I(AD15),
    .O(\BAR1/BR-15-8/RAWQ7 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND2   \BAR1/BR-15-8/$1I2960  (
    .I0(AD15),
    .I1(CFG53),
    .O(\BAR1/BR-15-8/IN7 )
  );
  X_AND2   \BAR1/BR-15-8/$1I2959  (
    .I0(CFG53),
    .I1(\BAR1/BR-15-8/RAWQ7 ),
    .O(\1BR15 )
  );
  X_AND2   \BAR1/BR-15-8/$1I2958  (
    .I0(CFG50),
    .I1(\BAR1/BR-15-8/RAWQ4 ),
    .O(\1BR12 )
  );
  X_AND2   \BAR1/BR-15-8/$1I2957  (
    .I0(CFG51),
    .I1(\BAR1/BR-15-8/RAWQ5 ),
    .O(\1BR13 )
  );
  X_AND2   \BAR1/BR-15-8/$1I2956  (
    .I0(AD13),
    .I1(CFG51),
    .O(\BAR1/BR-15-8/IN5 )
  );
  X_AND2   \BAR1/BR-15-8/$1I2955  (
    .I0(AD14),
    .I1(CFG52),
    .O(\BAR1/BR-15-8/IN6 )
  );
  X_AND2   \BAR1/BR-15-8/$1I2954  (
    .I0(CFG52),
    .I1(\BAR1/BR-15-8/RAWQ6 ),
    .O(\1BR14 )
  );
  X_XOR2   \BAR1/BR-15-8/X7  (
    .I0(\BAR1/BR-15-8/IN7 ),
    .I1(\1BR15 ),
    .O(\NlwInverterSignal_BAR1/BR-15-8/X7/O )
  );
  X_XOR2   \BAR1/BR-15-8/X5  (
    .I0(\BAR1/BR-15-8/IN5 ),
    .I1(\1BR13 ),
    .O(\NlwInverterSignal_BAR1/BR-15-8/X5/O )
  );
  X_ZERO   \BAR1/BR-15-8/$1I2909/$1I2218  (
    .O(\BAR1/BR-15-8/$1I2909/$1N2216 )
  );
  X_BUF   \BAR1/BR-15-8/$1I2909/L  (
    .I(\BAR1/BR-15-8/$1I2909/$1N2216 ),
    .O(\BAR1/BR-15-8/$1N2910 )
  );
  X_ZERO   \BAR1/BR-15-8/$1I2990/$1I2218  (
    .O(\BAR1/BR-15-8/$1I2990/$1N2216 )
  );
  X_BUF   \BAR1/BR-15-8/$1I2990/L  (
    .I(\BAR1/BR-15-8/$1I2990/$1N2216 ),
    .O(\BAR1/BR-15-8/$1N2911 )
  );
  X_ZERO   \BAR1/BR-15-8/$1I3091/$1I2218  (
    .O(\BAR1/BR-15-8/$1I3091/$1N2216 )
  );
  X_BUF   \BAR1/BR-15-8/$1I3091/L  (
    .I(\BAR1/BR-15-8/$1I3091/$1N2216 ),
    .O(\BAR1/BR-15-8/$1N3110 )
  );
  X_ZERO   \BAR1/BR-15-8/$1I3096/$1I2218  (
    .O(\BAR1/BR-15-8/$1I3096/$1N2216 )
  );
  X_BUF   \BAR1/BR-15-8/$1I3096/L  (
    .I(\BAR1/BR-15-8/$1I3096/$1N2216 ),
    .O(\BAR1/BR-15-8/$1N3111 )
  );
  X_INV   \BAR1/BR-CMD/$1I228  (
    .I(EX),
    .O(\BAR1/BR-CMD/EX_N )
  );
  X_AND3   \BAR1/BR-CMD/$1I194  (
    .I0(\NlwInverterSignal_BAR1/BR-CMD/$1I194/I0 ),
    .I1(CBE_IN3),
    .I2(CBE_IN2),
    .O(\BAR1/BR-CMD/$1N195 )
  );
  X_OR2   \BAR1/BR-CMD/$1I193  (
    .I0(\BAR1/BR-CMD/$1N195 ),
    .I1(\BAR1/BR-CMD/$1N201 ),
    .O(\BAR1/BR-CMD/MEM_6125 )
  );
  X_AND2   \BAR1/BR-CMD/$1I192  (
    .I0(CBE_IN2),
    .I1(CBE_IN1),
    .O(\BAR1/BR-CMD/$1N201 )
  );
  X_AND3   \BAR1/BR-CMD/$1I173  (
    .I0(\NlwInverterSignal_BAR1/BR-CMD/$1I173/I0 ),
    .I1(\NlwInverterSignal_BAR1/BR-CMD/$1I173/I1 ),
    .I2(CBE_IN1),
    .O(\BAR1/BR-CMD/IO_6122 )
  );
  X_MUX2   \BAR1/BR-CMD/$1I157  (
    .IB(\BAR1/$1N3380 ),
    .IA(\BAR1/BR-CMD/$1N144 ),
    .O(\BAR1/MATCH ),
    .SEL(\BAR1/BR-CMD/SEL )
  );
  X_AND2   \BAR1/BR-CMD/$1I117  (
    .I0(\NlwInverterSignal_BAR1/BR-CMD/$1I117/I0 ),
    .I1(CFG72),
    .O(\1BR2 )
  );
  X_AND2   \BAR1/BR-CMD/$1I110  (
    .I0(\NlwInverterSignal_BAR1/BR-CMD/$1I110/I0 ),
    .I1(CFG71),
    .O(\1BR1 )
  );
  X_BUF   \BAR1/BR-CMD/$1I109  (
    .I(CFG73),
    .O(\1BR0 )
  );
  X_AND2   \BAR1/BR-CMD/$1I100  (
    .I0(\NlwInverterSignal_BAR1/BR-CMD/$1I100/I0 ),
    .I1(CFG70),
    .O(\1BR3 )
  );
  X_ZERO   \BAR1/BR-CMD/$1I143/$1I2218  (
    .O(\BAR1/BR-CMD/$1I143/$1N2216 )
  );
  X_BUF   \BAR1/BR-CMD/$1I143/L  (
    .I(\BAR1/BR-CMD/$1I143/$1N2216 ),
    .O(\BAR1/BR-CMD/$1N144 )
  );
  X_OR2   \BAR1/BR-CMD/$1I223/$1I38  (
    .I0(\BAR1/BR-CMD/$1I223/M1 ),
    .I1(\BAR1/BR-CMD/$1I223/M0 ),
    .O(\BAR1/BR-CMD/SEL )
  );
  X_AND3   \BAR1/BR-CMD/$1I223/$1I31  (
    .I0(\NlwInverterSignal_BAR1/BR-CMD/$1I223/$1I31/I0 ),
    .I1(\BAR1/BR-CMD/EX_N ),
    .I2(\BAR1/BR-CMD/MEM_6125 ),
    .O(\BAR1/BR-CMD/$1I223/M0 )
  );
  X_AND3   \BAR1/BR-CMD/$1I223/$1I30  (
    .I0(\BAR1/BR-CMD/IO_6122 ),
    .I1(\BAR1/BR-CMD/EX_N ),
    .I2(CFG73),
    .O(\BAR1/BR-CMD/$1I223/M1 )
  );
  X_MUX2   \BAR1/BR-7-4/$1I2695  (
    .IB(CFG37),
    .IA(\BAR1/BR-7-4/$1N2701 ),
    .O(\BAR1/BR-7-4/$1N2697 ),
    .SEL(\BAR1/BR-7-4/EQ54_6161 )
  );
  X_MUX2   \BAR1/BR-7-4/$1I2694  (
    .IB(\BAR1/BR-7-4/$1N2697 ),
    .IA(\BAR1/BR-7-4/$1N2706 ),
    .O(\BAR1/$1N3366 ),
    .SEL(\BAR1/BR-7-4/EQ76_6160 )
  );
  X_AND2   \BAR1/BR-7-4/$1I2676  (
    .I0(AD4),
    .I1(CFG42),
    .O(\BAR1/BR-7-4/IN4 )
  );
  X_AND2   \BAR1/BR-7-4/$1I2672  (
    .I0(AD5),
    .I1(CFG43),
    .O(\BAR1/BR-7-4/IN5 )
  );
  X_AND2   \BAR1/BR-7-4/$1I2668  (
    .I0(AD6),
    .I1(CFG44),
    .O(\BAR1/BR-7-4/IN6 )
  );
  X_AND2   \BAR1/BR-7-4/$1I2664  (
    .I0(AD7),
    .I1(CFG45),
    .O(\BAR1/BR-7-4/IN7 )
  );
  X_AND2   \BAR1/BR-7-4/$1I2616  (
    .I0(CFG42),
    .I1(\BAR1/BR-7-4/RAWQ4 ),
    .O(\1BR4 )
  );
  X_AND2   \BAR1/BR-7-4/$1I2612  (
    .I0(CFG43),
    .I1(\BAR1/BR-7-4/RAWQ5 ),
    .O(\1BR5 )
  );
  X_AND2   \BAR1/BR-7-4/$1I2608  (
    .I0(CFG44),
    .I1(\BAR1/BR-7-4/RAWQ6 ),
    .O(\1BR6 )
  );
  X_AND2   \BAR1/BR-7-4/$1I2602  (
    .I0(CFG45),
    .I1(\BAR1/BR-7-4/RAWQ7 ),
    .O(\1BR7 )
  );
  X_AND2   \BAR1/BR-7-4/A2  (
    .I0(\BAR1/BR-7-4/EQ4 ),
    .I1(\BAR1/BR-7-4/EQ5 ),
    .O(\BAR1/BR-7-4/EQ54_6161 )
  );
  X_AND2   \BAR1/BR-7-4/A3  (
    .I0(\BAR1/BR-7-4/EQ6 ),
    .I1(\BAR1/BR-7-4/EQ7 ),
    .O(\BAR1/BR-7-4/EQ76_6160 )
  );
  X_XOR2   \BAR1/BR-7-4/X7  (
    .I0(\BAR1/BR-7-4/IN7 ),
    .I1(\1BR7 ),
    .O(\NlwInverterSignal_BAR1/BR-7-4/X7/O )
  );
  X_XOR2   \BAR1/BR-7-4/X6  (
    .I0(\BAR1/BR-7-4/IN6 ),
    .I1(\1BR6 ),
    .O(\NlwInverterSignal_BAR1/BR-7-4/X6/O )
  );
  X_XOR2   \BAR1/BR-7-4/X5  (
    .I0(\BAR1/BR-7-4/IN5 ),
    .I1(\1BR5 ),
    .O(\NlwInverterSignal_BAR1/BR-7-4/X5/O )
  );
  X_XOR2   \BAR1/BR-7-4/X4  (
    .I0(\BAR1/BR-7-4/IN4 ),
    .I1(\1BR4 ),
    .O(\NlwInverterSignal_BAR1/BR-7-4/X4/O )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR1/BR-7-4/Q7  (
    .CE(CE5_0),
    .CLK(CLK),
    .I(AD7),
    .O(\BAR1/BR-7-4/RAWQ7 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR1/BR-7-4/Q6  (
    .CE(CE5_0),
    .CLK(CLK),
    .I(AD6),
    .O(\BAR1/BR-7-4/RAWQ6 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR1/BR-7-4/Q5  (
    .CE(CE5_0),
    .CLK(CLK),
    .I(AD5),
    .O(\BAR1/BR-7-4/RAWQ5 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR1/BR-7-4/Q4  (
    .CE(CE5_0),
    .CLK(CLK),
    .I(AD4),
    .O(\BAR1/BR-7-4/RAWQ4 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_ZERO   \BAR1/BR-7-4/$1I2700/$1I2218  (
    .O(\BAR1/BR-7-4/$1I2700/$1N2216 )
  );
  X_BUF   \BAR1/BR-7-4/$1I2700/L  (
    .I(\BAR1/BR-7-4/$1I2700/$1N2216 ),
    .O(\BAR1/BR-7-4/$1N2701 )
  );
  X_ZERO   \BAR1/BR-7-4/$1I2705/$1I2218  (
    .O(\BAR1/BR-7-4/$1I2705/$1N2216 )
  );
  X_BUF   \BAR1/BR-7-4/$1I2705/L  (
    .I(\BAR1/BR-7-4/$1I2705/$1N2216 ),
    .O(\BAR1/BR-7-4/$1N2706 )
  );
  X_OR2   \BAR1/$1I3440/$1I38  (
    .I0(\BAR1/$1I3440/M1 ),
    .I1(\BAR1/$1I3440/M0 ),
    .O(\BAR1/CSREN32 )
  );
  X_AND3   \BAR1/$1I3440/$1I31  (
    .I0(\NlwInverterSignal_BAR1/$1I3440/$1I31/I0 ),
    .I1(CFG37),
    .I2(NlwRenamedSig_OI_CSR1),
    .O(\BAR1/$1I3440/M0 )
  );
  X_AND3   \BAR1/$1I3440/$1I30  (
    .I0(NlwRenamedSig_OI_CSR0),
    .I1(CFG37),
    .I2(CFG73),
    .O(\BAR1/$1I3440/M1 )
  );
  X_OR2   \BAR1/$1I3453/$1I38  (
    .I0(\BAR1/$1I3453/M1 ),
    .I1(\BAR1/$1I3453/M0 ),
    .O(\BAR1/CSREN64 )
  );
  X_AND3   \BAR1/$1I3453/$1I31  (
    .I0(\NlwInverterSignal_BAR1/$1I3453/$1I31/I0 ),
    .I1(CFG37),
    .I2(NlwRenamedSig_OI_CSR1),
    .O(\BAR1/$1I3453/M0 )
  );
  X_AND3   \BAR1/$1I3453/$1I30  (
    .I0(\BAR1/$1N3458 ),
    .I1(CFG37),
    .I2(CFG73),
    .O(\BAR1/$1I3453/M1 )
  );
  X_ZERO   \BAR1/$1I3468/$1I2218  (
    .O(\BAR1/$1I3468/$1N2216 )
  );
  X_BUF   \BAR1/$1I3468/L  (
    .I(\BAR1/$1I3468/$1N2216 ),
    .O(\BAR1/$1N3458 )
  );
  X_ONE   \BAR1/$1I3469/$1I2220  (
    .O(\BAR1/$1I3469/$1N2216 )
  );
  X_BUF   \BAR1/$1I3469/H  (
    .I(\BAR1/$1I3469/$1N2216 ),
    .O(\BAR1/ENABLE32 )
  );
  X_ONE   \BAR1/$2I3304/$1I2220  (
    .O(\BAR1/$2I3304/$1N2216 )
  );
  X_BUF   \BAR1/$2I3304/H  (
    .I(\BAR1/$2I3304/$1N2216 ),
    .O(\BAR1/ENABLENL )
  );
  X_OR2   \BAR1/$2I3321/$1I38  (
    .I0(\BAR1/$2I3321/M1 ),
    .I1(\BAR1/$2I3321/M0 ),
    .O(\BAR1/CSRENNL )
  );
  X_AND3   \BAR1/$2I3321/$1I31  (
    .I0(\NlwInverterSignal_BAR1/$2I3321/$1I31/I0 ),
    .I1(CFG37),
    .I2(NlwRenamedSig_OI_CSR1),
    .O(\BAR1/$2I3321/M0 )
  );
  X_AND3   \BAR1/$2I3321/$1I30  (
    .I0(NlwRenamedSig_OI_CSR0),
    .I1(CFG37),
    .I2(CFG73),
    .O(\BAR1/$2I3321/M1 )
  );
  X_AND4   \BAR2/$2I3324  (
    .I0(\BAR2/CSRENNL ),
    .I1(\BAR2/MATCH ),
    .I2(ADDR_VLD1),
    .I3(\BAR2/ENABLENL ),
    .O(\BAR2/NS_HITNL )
  );
  X_INV   \BAR2/$2I3284  (
    .I(CFG110),
    .O(\BAR2/NL_CE )
  );
  X_AND2   \BAR2/$2I3275  (
    .I0(\TSTOP_I- ),
    .I1(\BAR2/$2N3280 ),
    .O(\BAR2/NS_NL_MEM )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR2/NL  (
    .CE(\BAR2/NL_CE ),
    .CLK(CLK),
    .I(\BAR2/NS_NL_MEM ),
    .O(NL_MEM2),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_OR2   \BAR2/$2I3268  (
    .I0(\BAR2/$2N3273 ),
    .I1(NL_MEM2),
    .O(\BAR2/$2N3280 )
  );
  X_AND2   \BAR2/$2I3267  (
    .I0(\BAR2/UNALIGN ),
    .I1(\BAR2/NS_HITNL ),
    .O(\BAR2/$2N3273 )
  );
  X_OR2   \BAR2/$2I3263  (
    .I0(AD1),
    .I1(AD0),
    .O(\BAR2/UNALIGN )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR2/EQ64  (
    .CE(VCC),
    .CLK(CLK),
    .I(NS_BH64_2_INT),
    .O(BH64_2_INT),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR2/EQ32  (
    .CE(VCC),
    .CLK(CLK),
    .I(NS_BASE_HIT2_INT),
    .O(BASE_HIT2_INT),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND4   \BAR2/$1I3455  (
    .I0(\BAR2/CSREN64 ),
    .I1(\BAR2/MATCH ),
    .I2(ADDR_VLD64),
    .I3(CFG243),
    .O(NS_BH64_2_INT)
  );
  X_AND4   \BAR2/$1I3437  (
    .I0(\BAR2/CSREN32 ),
    .I1(\BAR2/MATCH ),
    .I2(ADDR_VLD1),
    .I3(\BAR2/ENABLE32 ),
    .O(NS_BASE_HIT2_INT)
  );
  X_MUX2   \BAR2/BR-31-24/$1I3094  (
    .IB(\BAR2/$1N3369 ),
    .IA(\BAR2/BR-31-24/$1N3110 ),
    .O(\BAR2/BR-31-24/$1N3099 ),
    .SEL(\BAR2/BR-31-24/EQ10_6397 )
  );
  X_MUX2   \BAR2/BR-31-24/$1I3093  (
    .IB(\BAR2/BR-31-24/$1N3099 ),
    .IA(\BAR2/BR-31-24/$1N3111 ),
    .O(\BAR2/BR-31-24/$1N2993 ),
    .SEL(\BAR2/BR-31-24/EQ32_6400 )
  );
  X_XOR2   \BAR2/BR-31-24/X1  (
    .I0(\BAR2/BR-31-24/IN1 ),
    .I1(\2BR25 ),
    .O(\NlwInverterSignal_BAR2/BR-31-24/X1/O )
  );
  X_XOR2   \BAR2/BR-31-24/X3  (
    .I0(\BAR2/BR-31-24/IN3 ),
    .I1(\2BR27 ),
    .O(\NlwInverterSignal_BAR2/BR-31-24/X3/O )
  );
  X_AND2   \BAR2/BR-31-24/$1I3014  (
    .I0(CFG101),
    .I1(\BAR2/BR-31-24/RAWQ2 ),
    .O(\2BR26 )
  );
  X_AND2   \BAR2/BR-31-24/$1I3013  (
    .I0(AD26),
    .I1(CFG101),
    .O(\BAR2/BR-31-24/IN2 )
  );
  X_AND2   \BAR2/BR-31-24/$1I3012  (
    .I0(AD25),
    .I1(CFG100),
    .O(\BAR2/BR-31-24/IN1 )
  );
  X_AND2   \BAR2/BR-31-24/$1I3011  (
    .I0(CFG100),
    .I1(\BAR2/BR-31-24/RAWQ1 ),
    .O(\2BR25 )
  );
  X_AND2   \BAR2/BR-31-24/$1I3010  (
    .I0(CFG99),
    .I1(\BAR2/BR-31-24/RAWQ0 ),
    .O(\2BR24 )
  );
  X_AND2   \BAR2/BR-31-24/$1I3009  (
    .I0(CFG102),
    .I1(\BAR2/BR-31-24/RAWQ3 ),
    .O(\2BR27 )
  );
  X_AND2   \BAR2/BR-31-24/$1I3008  (
    .I0(AD27),
    .I1(CFG102),
    .O(\BAR2/BR-31-24/IN3 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR2/BR-31-24/Q3  (
    .CE(CE6_3),
    .CLK(CLK),
    .I(AD27),
    .O(\BAR2/BR-31-24/RAWQ3 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR2/BR-31-24/Q2  (
    .CE(CE6_3),
    .CLK(CLK),
    .I(AD26),
    .O(\BAR2/BR-31-24/RAWQ2 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR2/BR-31-24/Q1  (
    .CE(CE6_3),
    .CLK(CLK),
    .I(AD25),
    .O(\BAR2/BR-31-24/RAWQ1 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR2/BR-31-24/Q0  (
    .CE(CE6_3),
    .CLK(CLK),
    .I(AD24),
    .O(\BAR2/BR-31-24/RAWQ0 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \BAR2/BR-31-24/X2  (
    .I0(\BAR2/BR-31-24/IN2 ),
    .I1(\2BR26 ),
    .O(\NlwInverterSignal_BAR2/BR-31-24/X2/O )
  );
  X_XOR2   \BAR2/BR-31-24/X0  (
    .I0(\BAR2/BR-31-24/IN0 ),
    .I1(\2BR24 ),
    .O(\NlwInverterSignal_BAR2/BR-31-24/X0/O )
  );
  X_AND2   \BAR2/BR-31-24/A1  (
    .I0(\BAR2/BR-31-24/EQ2 ),
    .I1(\BAR2/BR-31-24/EQ3 ),
    .O(\BAR2/BR-31-24/EQ32_6400 )
  );
  X_AND2   \BAR2/BR-31-24/A0  (
    .I0(\BAR2/BR-31-24/EQ0 ),
    .I1(\BAR2/BR-31-24/EQ1 ),
    .O(\BAR2/BR-31-24/EQ10_6397 )
  );
  X_AND2   \BAR2/BR-31-24/$1I2999  (
    .I0(AD24),
    .I1(CFG99),
    .O(\BAR2/BR-31-24/IN0 )
  );
  X_AND2   \BAR2/BR-31-24/$1I2989  (
    .I0(AD28),
    .I1(CFG103),
    .O(\BAR2/BR-31-24/IN4 )
  );
  X_AND2   \BAR2/BR-31-24/A2  (
    .I0(\BAR2/BR-31-24/EQ4 ),
    .I1(\BAR2/BR-31-24/EQ5 ),
    .O(\BAR2/BR-31-24/EQ54_6387 )
  );
  X_MUX2   \BAR2/BR-31-24/$1I2986  (
    .IB(\BAR2/BR-31-24/$1N2992 ),
    .IA(\BAR2/BR-31-24/$1N2910 ),
    .O(\BAR2/$1N3380 ),
    .SEL(\BAR2/BR-31-24/EQ76_6390 )
  );
  X_MUX2   \BAR2/BR-31-24/$1I2985  (
    .IB(\BAR2/BR-31-24/$1N2993 ),
    .IA(\BAR2/BR-31-24/$1N2911 ),
    .O(\BAR2/BR-31-24/$1N2992 ),
    .SEL(\BAR2/BR-31-24/EQ54_6387 )
  );
  X_AND2   \BAR2/BR-31-24/A3  (
    .I0(\BAR2/BR-31-24/EQ6 ),
    .I1(\BAR2/BR-31-24/EQ7 ),
    .O(\BAR2/BR-31-24/EQ76_6390 )
  );
  X_XOR2   \BAR2/BR-31-24/X4  (
    .I0(\BAR2/BR-31-24/IN4 ),
    .I1(\2BR28 ),
    .O(\NlwInverterSignal_BAR2/BR-31-24/X4/O )
  );
  X_XOR2   \BAR2/BR-31-24/X6  (
    .I0(\BAR2/BR-31-24/IN6 ),
    .I1(\2BR30 ),
    .O(\NlwInverterSignal_BAR2/BR-31-24/X6/O )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR2/BR-31-24/Q4  (
    .CE(CE6_3),
    .CLK(CLK),
    .I(AD28),
    .O(\BAR2/BR-31-24/RAWQ4 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR2/BR-31-24/Q5  (
    .CE(CE6_3),
    .CLK(CLK),
    .I(AD29),
    .O(\BAR2/BR-31-24/RAWQ5 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR2/BR-31-24/Q6  (
    .CE(CE6_3),
    .CLK(CLK),
    .I(AD30),
    .O(\BAR2/BR-31-24/RAWQ6 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR2/BR-31-24/Q7  (
    .CE(CE6_3),
    .CLK(CLK),
    .I(AD31),
    .O(\BAR2/BR-31-24/RAWQ7 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND2   \BAR2/BR-31-24/$1I2960  (
    .I0(AD31),
    .I1(CFG106),
    .O(\BAR2/BR-31-24/IN7 )
  );
  X_AND2   \BAR2/BR-31-24/$1I2959  (
    .I0(CFG106),
    .I1(\BAR2/BR-31-24/RAWQ7 ),
    .O(\2BR31 )
  );
  X_AND2   \BAR2/BR-31-24/$1I2958  (
    .I0(CFG103),
    .I1(\BAR2/BR-31-24/RAWQ4 ),
    .O(\2BR28 )
  );
  X_AND2   \BAR2/BR-31-24/$1I2957  (
    .I0(CFG104),
    .I1(\BAR2/BR-31-24/RAWQ5 ),
    .O(\2BR29 )
  );
  X_AND2   \BAR2/BR-31-24/$1I2956  (
    .I0(AD29),
    .I1(CFG104),
    .O(\BAR2/BR-31-24/IN5 )
  );
  X_AND2   \BAR2/BR-31-24/$1I2955  (
    .I0(AD30),
    .I1(CFG105),
    .O(\BAR2/BR-31-24/IN6 )
  );
  X_AND2   \BAR2/BR-31-24/$1I2954  (
    .I0(CFG105),
    .I1(\BAR2/BR-31-24/RAWQ6 ),
    .O(\2BR30 )
  );
  X_XOR2   \BAR2/BR-31-24/X7  (
    .I0(\BAR2/BR-31-24/IN7 ),
    .I1(\2BR31 ),
    .O(\NlwInverterSignal_BAR2/BR-31-24/X7/O )
  );
  X_XOR2   \BAR2/BR-31-24/X5  (
    .I0(\BAR2/BR-31-24/IN5 ),
    .I1(\2BR29 ),
    .O(\NlwInverterSignal_BAR2/BR-31-24/X5/O )
  );
  X_ZERO   \BAR2/BR-31-24/$1I2909/$1I2218  (
    .O(\BAR2/BR-31-24/$1I2909/$1N2216 )
  );
  X_BUF   \BAR2/BR-31-24/$1I2909/L  (
    .I(\BAR2/BR-31-24/$1I2909/$1N2216 ),
    .O(\BAR2/BR-31-24/$1N2910 )
  );
  X_ZERO   \BAR2/BR-31-24/$1I2990/$1I2218  (
    .O(\BAR2/BR-31-24/$1I2990/$1N2216 )
  );
  X_BUF   \BAR2/BR-31-24/$1I2990/L  (
    .I(\BAR2/BR-31-24/$1I2990/$1N2216 ),
    .O(\BAR2/BR-31-24/$1N2911 )
  );
  X_ZERO   \BAR2/BR-31-24/$1I3091/$1I2218  (
    .O(\BAR2/BR-31-24/$1I3091/$1N2216 )
  );
  X_BUF   \BAR2/BR-31-24/$1I3091/L  (
    .I(\BAR2/BR-31-24/$1I3091/$1N2216 ),
    .O(\BAR2/BR-31-24/$1N3110 )
  );
  X_ZERO   \BAR2/BR-31-24/$1I3096/$1I2218  (
    .O(\BAR2/BR-31-24/$1I3096/$1N2216 )
  );
  X_BUF   \BAR2/BR-31-24/$1I3096/L  (
    .I(\BAR2/BR-31-24/$1I3096/$1N2216 ),
    .O(\BAR2/BR-31-24/$1N3111 )
  );
  X_MUX2   \BAR2/BR-23-16/$1I3094  (
    .IB(\BAR2/$1N3368 ),
    .IA(\BAR2/BR-23-16/$1N3110 ),
    .O(\BAR2/BR-23-16/$1N3099 ),
    .SEL(\BAR2/BR-23-16/EQ10_6469 )
  );
  X_MUX2   \BAR2/BR-23-16/$1I3093  (
    .IB(\BAR2/BR-23-16/$1N3099 ),
    .IA(\BAR2/BR-23-16/$1N3111 ),
    .O(\BAR2/BR-23-16/$1N2993 ),
    .SEL(\BAR2/BR-23-16/EQ32_6472 )
  );
  X_XOR2   \BAR2/BR-23-16/X1  (
    .I0(\BAR2/BR-23-16/IN1 ),
    .I1(\2BR17 ),
    .O(\NlwInverterSignal_BAR2/BR-23-16/X1/O )
  );
  X_XOR2   \BAR2/BR-23-16/X3  (
    .I0(\BAR2/BR-23-16/IN3 ),
    .I1(\2BR19 ),
    .O(\NlwInverterSignal_BAR2/BR-23-16/X3/O )
  );
  X_AND2   \BAR2/BR-23-16/$1I3014  (
    .I0(CFG93),
    .I1(\BAR2/BR-23-16/RAWQ2 ),
    .O(\2BR18 )
  );
  X_AND2   \BAR2/BR-23-16/$1I3013  (
    .I0(AD18),
    .I1(CFG93),
    .O(\BAR2/BR-23-16/IN2 )
  );
  X_AND2   \BAR2/BR-23-16/$1I3012  (
    .I0(AD17),
    .I1(CFG92),
    .O(\BAR2/BR-23-16/IN1 )
  );
  X_AND2   \BAR2/BR-23-16/$1I3011  (
    .I0(CFG92),
    .I1(\BAR2/BR-23-16/RAWQ1 ),
    .O(\2BR17 )
  );
  X_AND2   \BAR2/BR-23-16/$1I3010  (
    .I0(CFG91),
    .I1(\BAR2/BR-23-16/RAWQ0 ),
    .O(\2BR16 )
  );
  X_AND2   \BAR2/BR-23-16/$1I3009  (
    .I0(CFG94),
    .I1(\BAR2/BR-23-16/RAWQ3 ),
    .O(\2BR19 )
  );
  X_AND2   \BAR2/BR-23-16/$1I3008  (
    .I0(AD19),
    .I1(CFG94),
    .O(\BAR2/BR-23-16/IN3 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR2/BR-23-16/Q3  (
    .CE(CE6_2),
    .CLK(CLK),
    .I(AD19),
    .O(\BAR2/BR-23-16/RAWQ3 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR2/BR-23-16/Q2  (
    .CE(CE6_2),
    .CLK(CLK),
    .I(AD18),
    .O(\BAR2/BR-23-16/RAWQ2 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR2/BR-23-16/Q1  (
    .CE(CE6_2),
    .CLK(CLK),
    .I(AD17),
    .O(\BAR2/BR-23-16/RAWQ1 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR2/BR-23-16/Q0  (
    .CE(CE6_2),
    .CLK(CLK),
    .I(AD16),
    .O(\BAR2/BR-23-16/RAWQ0 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \BAR2/BR-23-16/X2  (
    .I0(\BAR2/BR-23-16/IN2 ),
    .I1(\2BR18 ),
    .O(\NlwInverterSignal_BAR2/BR-23-16/X2/O )
  );
  X_XOR2   \BAR2/BR-23-16/X0  (
    .I0(\BAR2/BR-23-16/IN0 ),
    .I1(\2BR16 ),
    .O(\NlwInverterSignal_BAR2/BR-23-16/X0/O )
  );
  X_AND2   \BAR2/BR-23-16/A1  (
    .I0(\BAR2/BR-23-16/EQ2 ),
    .I1(\BAR2/BR-23-16/EQ3 ),
    .O(\BAR2/BR-23-16/EQ32_6472 )
  );
  X_AND2   \BAR2/BR-23-16/A0  (
    .I0(\BAR2/BR-23-16/EQ0 ),
    .I1(\BAR2/BR-23-16/EQ1 ),
    .O(\BAR2/BR-23-16/EQ10_6469 )
  );
  X_AND2   \BAR2/BR-23-16/$1I2999  (
    .I0(AD16),
    .I1(CFG91),
    .O(\BAR2/BR-23-16/IN0 )
  );
  X_AND2   \BAR2/BR-23-16/$1I2989  (
    .I0(AD20),
    .I1(CFG95),
    .O(\BAR2/BR-23-16/IN4 )
  );
  X_AND2   \BAR2/BR-23-16/A2  (
    .I0(\BAR2/BR-23-16/EQ4 ),
    .I1(\BAR2/BR-23-16/EQ5 ),
    .O(\BAR2/BR-23-16/EQ54_6459 )
  );
  X_MUX2   \BAR2/BR-23-16/$1I2986  (
    .IB(\BAR2/BR-23-16/$1N2992 ),
    .IA(\BAR2/BR-23-16/$1N2910 ),
    .O(\BAR2/$1N3369 ),
    .SEL(\BAR2/BR-23-16/EQ76_6462 )
  );
  X_MUX2   \BAR2/BR-23-16/$1I2985  (
    .IB(\BAR2/BR-23-16/$1N2993 ),
    .IA(\BAR2/BR-23-16/$1N2911 ),
    .O(\BAR2/BR-23-16/$1N2992 ),
    .SEL(\BAR2/BR-23-16/EQ54_6459 )
  );
  X_AND2   \BAR2/BR-23-16/A3  (
    .I0(\BAR2/BR-23-16/EQ6 ),
    .I1(\BAR2/BR-23-16/EQ7 ),
    .O(\BAR2/BR-23-16/EQ76_6462 )
  );
  X_XOR2   \BAR2/BR-23-16/X4  (
    .I0(\BAR2/BR-23-16/IN4 ),
    .I1(\2BR20 ),
    .O(\NlwInverterSignal_BAR2/BR-23-16/X4/O )
  );
  X_XOR2   \BAR2/BR-23-16/X6  (
    .I0(\BAR2/BR-23-16/IN6 ),
    .I1(\2BR22 ),
    .O(\NlwInverterSignal_BAR2/BR-23-16/X6/O )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR2/BR-23-16/Q4  (
    .CE(CE6_2),
    .CLK(CLK),
    .I(AD20),
    .O(\BAR2/BR-23-16/RAWQ4 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR2/BR-23-16/Q5  (
    .CE(CE6_2),
    .CLK(CLK),
    .I(AD21),
    .O(\BAR2/BR-23-16/RAWQ5 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR2/BR-23-16/Q6  (
    .CE(CE6_2),
    .CLK(CLK),
    .I(AD22),
    .O(\BAR2/BR-23-16/RAWQ6 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR2/BR-23-16/Q7  (
    .CE(CE6_2),
    .CLK(CLK),
    .I(AD23),
    .O(\BAR2/BR-23-16/RAWQ7 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND2   \BAR2/BR-23-16/$1I2960  (
    .I0(AD23),
    .I1(CFG98),
    .O(\BAR2/BR-23-16/IN7 )
  );
  X_AND2   \BAR2/BR-23-16/$1I2959  (
    .I0(CFG98),
    .I1(\BAR2/BR-23-16/RAWQ7 ),
    .O(\2BR23 )
  );
  X_AND2   \BAR2/BR-23-16/$1I2958  (
    .I0(CFG95),
    .I1(\BAR2/BR-23-16/RAWQ4 ),
    .O(\2BR20 )
  );
  X_AND2   \BAR2/BR-23-16/$1I2957  (
    .I0(CFG96),
    .I1(\BAR2/BR-23-16/RAWQ5 ),
    .O(\2BR21 )
  );
  X_AND2   \BAR2/BR-23-16/$1I2956  (
    .I0(AD21),
    .I1(CFG96),
    .O(\BAR2/BR-23-16/IN5 )
  );
  X_AND2   \BAR2/BR-23-16/$1I2955  (
    .I0(AD22),
    .I1(CFG97),
    .O(\BAR2/BR-23-16/IN6 )
  );
  X_AND2   \BAR2/BR-23-16/$1I2954  (
    .I0(CFG97),
    .I1(\BAR2/BR-23-16/RAWQ6 ),
    .O(\2BR22 )
  );
  X_XOR2   \BAR2/BR-23-16/X7  (
    .I0(\BAR2/BR-23-16/IN7 ),
    .I1(\2BR23 ),
    .O(\NlwInverterSignal_BAR2/BR-23-16/X7/O )
  );
  X_XOR2   \BAR2/BR-23-16/X5  (
    .I0(\BAR2/BR-23-16/IN5 ),
    .I1(\2BR21 ),
    .O(\NlwInverterSignal_BAR2/BR-23-16/X5/O )
  );
  X_ZERO   \BAR2/BR-23-16/$1I2909/$1I2218  (
    .O(\BAR2/BR-23-16/$1I2909/$1N2216 )
  );
  X_BUF   \BAR2/BR-23-16/$1I2909/L  (
    .I(\BAR2/BR-23-16/$1I2909/$1N2216 ),
    .O(\BAR2/BR-23-16/$1N2910 )
  );
  X_ZERO   \BAR2/BR-23-16/$1I2990/$1I2218  (
    .O(\BAR2/BR-23-16/$1I2990/$1N2216 )
  );
  X_BUF   \BAR2/BR-23-16/$1I2990/L  (
    .I(\BAR2/BR-23-16/$1I2990/$1N2216 ),
    .O(\BAR2/BR-23-16/$1N2911 )
  );
  X_ZERO   \BAR2/BR-23-16/$1I3091/$1I2218  (
    .O(\BAR2/BR-23-16/$1I3091/$1N2216 )
  );
  X_BUF   \BAR2/BR-23-16/$1I3091/L  (
    .I(\BAR2/BR-23-16/$1I3091/$1N2216 ),
    .O(\BAR2/BR-23-16/$1N3110 )
  );
  X_ZERO   \BAR2/BR-23-16/$1I3096/$1I2218  (
    .O(\BAR2/BR-23-16/$1I3096/$1N2216 )
  );
  X_BUF   \BAR2/BR-23-16/$1I3096/L  (
    .I(\BAR2/BR-23-16/$1I3096/$1N2216 ),
    .O(\BAR2/BR-23-16/$1N3111 )
  );
  X_MUX2   \BAR2/BR-15-8/$1I3094  (
    .IB(\BAR2/$1N3366 ),
    .IA(\BAR2/BR-15-8/$1N3110 ),
    .O(\BAR2/BR-15-8/$1N3099 ),
    .SEL(\BAR2/BR-15-8/EQ10_6541 )
  );
  X_MUX2   \BAR2/BR-15-8/$1I3093  (
    .IB(\BAR2/BR-15-8/$1N3099 ),
    .IA(\BAR2/BR-15-8/$1N3111 ),
    .O(\BAR2/BR-15-8/$1N2993 ),
    .SEL(\BAR2/BR-15-8/EQ32_6544 )
  );
  X_XOR2   \BAR2/BR-15-8/X1  (
    .I0(\BAR2/BR-15-8/IN1 ),
    .I1(\2BR9 ),
    .O(\NlwInverterSignal_BAR2/BR-15-8/X1/O )
  );
  X_XOR2   \BAR2/BR-15-8/X3  (
    .I0(\BAR2/BR-15-8/IN3 ),
    .I1(\2BR11 ),
    .O(\NlwInverterSignal_BAR2/BR-15-8/X3/O )
  );
  X_AND2   \BAR2/BR-15-8/$1I3014  (
    .I0(CFG85),
    .I1(\BAR2/BR-15-8/RAWQ2 ),
    .O(\2BR10 )
  );
  X_AND2   \BAR2/BR-15-8/$1I3013  (
    .I0(AD10),
    .I1(CFG85),
    .O(\BAR2/BR-15-8/IN2 )
  );
  X_AND2   \BAR2/BR-15-8/$1I3012  (
    .I0(AD9),
    .I1(CFG84),
    .O(\BAR2/BR-15-8/IN1 )
  );
  X_AND2   \BAR2/BR-15-8/$1I3011  (
    .I0(CFG84),
    .I1(\BAR2/BR-15-8/RAWQ1 ),
    .O(\2BR9 )
  );
  X_AND2   \BAR2/BR-15-8/$1I3010  (
    .I0(CFG83),
    .I1(\BAR2/BR-15-8/RAWQ0 ),
    .O(\2BR8 )
  );
  X_AND2   \BAR2/BR-15-8/$1I3009  (
    .I0(CFG86),
    .I1(\BAR2/BR-15-8/RAWQ3 ),
    .O(\2BR11 )
  );
  X_AND2   \BAR2/BR-15-8/$1I3008  (
    .I0(AD11),
    .I1(CFG86),
    .O(\BAR2/BR-15-8/IN3 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR2/BR-15-8/Q3  (
    .CE(CE6_1),
    .CLK(CLK),
    .I(AD11),
    .O(\BAR2/BR-15-8/RAWQ3 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR2/BR-15-8/Q2  (
    .CE(CE6_1),
    .CLK(CLK),
    .I(AD10),
    .O(\BAR2/BR-15-8/RAWQ2 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR2/BR-15-8/Q1  (
    .CE(CE6_1),
    .CLK(CLK),
    .I(AD9),
    .O(\BAR2/BR-15-8/RAWQ1 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR2/BR-15-8/Q0  (
    .CE(CE6_1),
    .CLK(CLK),
    .I(AD8),
    .O(\BAR2/BR-15-8/RAWQ0 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \BAR2/BR-15-8/X2  (
    .I0(\BAR2/BR-15-8/IN2 ),
    .I1(\2BR10 ),
    .O(\NlwInverterSignal_BAR2/BR-15-8/X2/O )
  );
  X_XOR2   \BAR2/BR-15-8/X0  (
    .I0(\BAR2/BR-15-8/IN0 ),
    .I1(\2BR8 ),
    .O(\NlwInverterSignal_BAR2/BR-15-8/X0/O )
  );
  X_AND2   \BAR2/BR-15-8/A1  (
    .I0(\BAR2/BR-15-8/EQ2 ),
    .I1(\BAR2/BR-15-8/EQ3 ),
    .O(\BAR2/BR-15-8/EQ32_6544 )
  );
  X_AND2   \BAR2/BR-15-8/A0  (
    .I0(\BAR2/BR-15-8/EQ0 ),
    .I1(\BAR2/BR-15-8/EQ1 ),
    .O(\BAR2/BR-15-8/EQ10_6541 )
  );
  X_AND2   \BAR2/BR-15-8/$1I2999  (
    .I0(AD8),
    .I1(CFG83),
    .O(\BAR2/BR-15-8/IN0 )
  );
  X_AND2   \BAR2/BR-15-8/$1I2989  (
    .I0(AD12),
    .I1(CFG87),
    .O(\BAR2/BR-15-8/IN4 )
  );
  X_AND2   \BAR2/BR-15-8/A2  (
    .I0(\BAR2/BR-15-8/EQ4 ),
    .I1(\BAR2/BR-15-8/EQ5 ),
    .O(\BAR2/BR-15-8/EQ54_6531 )
  );
  X_MUX2   \BAR2/BR-15-8/$1I2986  (
    .IB(\BAR2/BR-15-8/$1N2992 ),
    .IA(\BAR2/BR-15-8/$1N2910 ),
    .O(\BAR2/$1N3368 ),
    .SEL(\BAR2/BR-15-8/EQ76_6534 )
  );
  X_MUX2   \BAR2/BR-15-8/$1I2985  (
    .IB(\BAR2/BR-15-8/$1N2993 ),
    .IA(\BAR2/BR-15-8/$1N2911 ),
    .O(\BAR2/BR-15-8/$1N2992 ),
    .SEL(\BAR2/BR-15-8/EQ54_6531 )
  );
  X_AND2   \BAR2/BR-15-8/A3  (
    .I0(\BAR2/BR-15-8/EQ6 ),
    .I1(\BAR2/BR-15-8/EQ7 ),
    .O(\BAR2/BR-15-8/EQ76_6534 )
  );
  X_XOR2   \BAR2/BR-15-8/X4  (
    .I0(\BAR2/BR-15-8/IN4 ),
    .I1(\2BR12 ),
    .O(\NlwInverterSignal_BAR2/BR-15-8/X4/O )
  );
  X_XOR2   \BAR2/BR-15-8/X6  (
    .I0(\BAR2/BR-15-8/IN6 ),
    .I1(\2BR14 ),
    .O(\NlwInverterSignal_BAR2/BR-15-8/X6/O )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR2/BR-15-8/Q4  (
    .CE(CE6_1),
    .CLK(CLK),
    .I(AD12),
    .O(\BAR2/BR-15-8/RAWQ4 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR2/BR-15-8/Q5  (
    .CE(CE6_1),
    .CLK(CLK),
    .I(AD13),
    .O(\BAR2/BR-15-8/RAWQ5 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR2/BR-15-8/Q6  (
    .CE(CE6_1),
    .CLK(CLK),
    .I(AD14),
    .O(\BAR2/BR-15-8/RAWQ6 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR2/BR-15-8/Q7  (
    .CE(CE6_1),
    .CLK(CLK),
    .I(AD15),
    .O(\BAR2/BR-15-8/RAWQ7 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND2   \BAR2/BR-15-8/$1I2960  (
    .I0(AD15),
    .I1(CFG90),
    .O(\BAR2/BR-15-8/IN7 )
  );
  X_AND2   \BAR2/BR-15-8/$1I2959  (
    .I0(CFG90),
    .I1(\BAR2/BR-15-8/RAWQ7 ),
    .O(\2BR15 )
  );
  X_AND2   \BAR2/BR-15-8/$1I2958  (
    .I0(CFG87),
    .I1(\BAR2/BR-15-8/RAWQ4 ),
    .O(\2BR12 )
  );
  X_AND2   \BAR2/BR-15-8/$1I2957  (
    .I0(CFG88),
    .I1(\BAR2/BR-15-8/RAWQ5 ),
    .O(\2BR13 )
  );
  X_AND2   \BAR2/BR-15-8/$1I2956  (
    .I0(AD13),
    .I1(CFG88),
    .O(\BAR2/BR-15-8/IN5 )
  );
  X_AND2   \BAR2/BR-15-8/$1I2955  (
    .I0(AD14),
    .I1(CFG89),
    .O(\BAR2/BR-15-8/IN6 )
  );
  X_AND2   \BAR2/BR-15-8/$1I2954  (
    .I0(CFG89),
    .I1(\BAR2/BR-15-8/RAWQ6 ),
    .O(\2BR14 )
  );
  X_XOR2   \BAR2/BR-15-8/X7  (
    .I0(\BAR2/BR-15-8/IN7 ),
    .I1(\2BR15 ),
    .O(\NlwInverterSignal_BAR2/BR-15-8/X7/O )
  );
  X_XOR2   \BAR2/BR-15-8/X5  (
    .I0(\BAR2/BR-15-8/IN5 ),
    .I1(\2BR13 ),
    .O(\NlwInverterSignal_BAR2/BR-15-8/X5/O )
  );
  X_ZERO   \BAR2/BR-15-8/$1I2909/$1I2218  (
    .O(\BAR2/BR-15-8/$1I2909/$1N2216 )
  );
  X_BUF   \BAR2/BR-15-8/$1I2909/L  (
    .I(\BAR2/BR-15-8/$1I2909/$1N2216 ),
    .O(\BAR2/BR-15-8/$1N2910 )
  );
  X_ZERO   \BAR2/BR-15-8/$1I2990/$1I2218  (
    .O(\BAR2/BR-15-8/$1I2990/$1N2216 )
  );
  X_BUF   \BAR2/BR-15-8/$1I2990/L  (
    .I(\BAR2/BR-15-8/$1I2990/$1N2216 ),
    .O(\BAR2/BR-15-8/$1N2911 )
  );
  X_ZERO   \BAR2/BR-15-8/$1I3091/$1I2218  (
    .O(\BAR2/BR-15-8/$1I3091/$1N2216 )
  );
  X_BUF   \BAR2/BR-15-8/$1I3091/L  (
    .I(\BAR2/BR-15-8/$1I3091/$1N2216 ),
    .O(\BAR2/BR-15-8/$1N3110 )
  );
  X_ZERO   \BAR2/BR-15-8/$1I3096/$1I2218  (
    .O(\BAR2/BR-15-8/$1I3096/$1N2216 )
  );
  X_BUF   \BAR2/BR-15-8/$1I3096/L  (
    .I(\BAR2/BR-15-8/$1I3096/$1N2216 ),
    .O(\BAR2/BR-15-8/$1N3111 )
  );
  X_INV   \BAR2/BR-CMD/$1I228  (
    .I(EX),
    .O(\BAR2/BR-CMD/EX_N )
  );
  X_AND3   \BAR2/BR-CMD/$1I194  (
    .I0(\NlwInverterSignal_BAR2/BR-CMD/$1I194/I0 ),
    .I1(CBE_IN3),
    .I2(CBE_IN2),
    .O(\BAR2/BR-CMD/$1N195 )
  );
  X_OR2   \BAR2/BR-CMD/$1I193  (
    .I0(\BAR2/BR-CMD/$1N195 ),
    .I1(\BAR2/BR-CMD/$1N201 ),
    .O(\BAR2/BR-CMD/MEM_6584 )
  );
  X_AND2   \BAR2/BR-CMD/$1I192  (
    .I0(CBE_IN2),
    .I1(CBE_IN1),
    .O(\BAR2/BR-CMD/$1N201 )
  );
  X_AND3   \BAR2/BR-CMD/$1I173  (
    .I0(\NlwInverterSignal_BAR2/BR-CMD/$1I173/I0 ),
    .I1(\NlwInverterSignal_BAR2/BR-CMD/$1I173/I1 ),
    .I2(CBE_IN1),
    .O(\BAR2/BR-CMD/IO_6581 )
  );
  X_MUX2   \BAR2/BR-CMD/$1I157  (
    .IB(\BAR2/$1N3380 ),
    .IA(\BAR2/BR-CMD/$1N144 ),
    .O(\BAR2/MATCH ),
    .SEL(\BAR2/BR-CMD/SEL )
  );
  X_AND2   \BAR2/BR-CMD/$1I117  (
    .I0(\NlwInverterSignal_BAR2/BR-CMD/$1I117/I0 ),
    .I1(CFG109),
    .O(\2BR2 )
  );
  X_AND2   \BAR2/BR-CMD/$1I110  (
    .I0(\NlwInverterSignal_BAR2/BR-CMD/$1I110/I0 ),
    .I1(CFG108),
    .O(\2BR1 )
  );
  X_BUF   \BAR2/BR-CMD/$1I109  (
    .I(CFG110),
    .O(\2BR0 )
  );
  X_AND2   \BAR2/BR-CMD/$1I100  (
    .I0(\NlwInverterSignal_BAR2/BR-CMD/$1I100/I0 ),
    .I1(CFG107),
    .O(\2BR3 )
  );
  X_ZERO   \BAR2/BR-CMD/$1I143/$1I2218  (
    .O(\BAR2/BR-CMD/$1I143/$1N2216 )
  );
  X_BUF   \BAR2/BR-CMD/$1I143/L  (
    .I(\BAR2/BR-CMD/$1I143/$1N2216 ),
    .O(\BAR2/BR-CMD/$1N144 )
  );
  X_OR2   \BAR2/BR-CMD/$1I223/$1I38  (
    .I0(\BAR2/BR-CMD/$1I223/M1 ),
    .I1(\BAR2/BR-CMD/$1I223/M0 ),
    .O(\BAR2/BR-CMD/SEL )
  );
  X_AND3   \BAR2/BR-CMD/$1I223/$1I31  (
    .I0(\NlwInverterSignal_BAR2/BR-CMD/$1I223/$1I31/I0 ),
    .I1(\BAR2/BR-CMD/EX_N ),
    .I2(\BAR2/BR-CMD/MEM_6584 ),
    .O(\BAR2/BR-CMD/$1I223/M0 )
  );
  X_AND3   \BAR2/BR-CMD/$1I223/$1I30  (
    .I0(\BAR2/BR-CMD/IO_6581 ),
    .I1(\BAR2/BR-CMD/EX_N ),
    .I2(CFG110),
    .O(\BAR2/BR-CMD/$1I223/M1 )
  );
  X_MUX2   \BAR2/BR-7-4/$1I2695  (
    .IB(CFG74),
    .IA(\BAR2/BR-7-4/$1N2701 ),
    .O(\BAR2/BR-7-4/$1N2697 ),
    .SEL(\BAR2/BR-7-4/EQ54_6620 )
  );
  X_MUX2   \BAR2/BR-7-4/$1I2694  (
    .IB(\BAR2/BR-7-4/$1N2697 ),
    .IA(\BAR2/BR-7-4/$1N2706 ),
    .O(\BAR2/$1N3366 ),
    .SEL(\BAR2/BR-7-4/EQ76_6619 )
  );
  X_AND2   \BAR2/BR-7-4/$1I2676  (
    .I0(AD4),
    .I1(CFG79),
    .O(\BAR2/BR-7-4/IN4 )
  );
  X_AND2   \BAR2/BR-7-4/$1I2672  (
    .I0(AD5),
    .I1(CFG80),
    .O(\BAR2/BR-7-4/IN5 )
  );
  X_AND2   \BAR2/BR-7-4/$1I2668  (
    .I0(AD6),
    .I1(CFG81),
    .O(\BAR2/BR-7-4/IN6 )
  );
  X_AND2   \BAR2/BR-7-4/$1I2664  (
    .I0(AD7),
    .I1(CFG82),
    .O(\BAR2/BR-7-4/IN7 )
  );
  X_AND2   \BAR2/BR-7-4/$1I2616  (
    .I0(CFG79),
    .I1(\BAR2/BR-7-4/RAWQ4 ),
    .O(\2BR4 )
  );
  X_AND2   \BAR2/BR-7-4/$1I2612  (
    .I0(CFG80),
    .I1(\BAR2/BR-7-4/RAWQ5 ),
    .O(\2BR5 )
  );
  X_AND2   \BAR2/BR-7-4/$1I2608  (
    .I0(CFG81),
    .I1(\BAR2/BR-7-4/RAWQ6 ),
    .O(\2BR6 )
  );
  X_AND2   \BAR2/BR-7-4/$1I2602  (
    .I0(CFG82),
    .I1(\BAR2/BR-7-4/RAWQ7 ),
    .O(\2BR7 )
  );
  X_AND2   \BAR2/BR-7-4/A2  (
    .I0(\BAR2/BR-7-4/EQ4 ),
    .I1(\BAR2/BR-7-4/EQ5 ),
    .O(\BAR2/BR-7-4/EQ54_6620 )
  );
  X_AND2   \BAR2/BR-7-4/A3  (
    .I0(\BAR2/BR-7-4/EQ6 ),
    .I1(\BAR2/BR-7-4/EQ7 ),
    .O(\BAR2/BR-7-4/EQ76_6619 )
  );
  X_XOR2   \BAR2/BR-7-4/X7  (
    .I0(\BAR2/BR-7-4/IN7 ),
    .I1(\2BR7 ),
    .O(\NlwInverterSignal_BAR2/BR-7-4/X7/O )
  );
  X_XOR2   \BAR2/BR-7-4/X6  (
    .I0(\BAR2/BR-7-4/IN6 ),
    .I1(\2BR6 ),
    .O(\NlwInverterSignal_BAR2/BR-7-4/X6/O )
  );
  X_XOR2   \BAR2/BR-7-4/X5  (
    .I0(\BAR2/BR-7-4/IN5 ),
    .I1(\2BR5 ),
    .O(\NlwInverterSignal_BAR2/BR-7-4/X5/O )
  );
  X_XOR2   \BAR2/BR-7-4/X4  (
    .I0(\BAR2/BR-7-4/IN4 ),
    .I1(\2BR4 ),
    .O(\NlwInverterSignal_BAR2/BR-7-4/X4/O )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR2/BR-7-4/Q7  (
    .CE(CE6_0),
    .CLK(CLK),
    .I(AD7),
    .O(\BAR2/BR-7-4/RAWQ7 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR2/BR-7-4/Q6  (
    .CE(CE6_0),
    .CLK(CLK),
    .I(AD6),
    .O(\BAR2/BR-7-4/RAWQ6 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR2/BR-7-4/Q5  (
    .CE(CE6_0),
    .CLK(CLK),
    .I(AD5),
    .O(\BAR2/BR-7-4/RAWQ5 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \BAR2/BR-7-4/Q4  (
    .CE(CE6_0),
    .CLK(CLK),
    .I(AD4),
    .O(\BAR2/BR-7-4/RAWQ4 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_ZERO   \BAR2/BR-7-4/$1I2700/$1I2218  (
    .O(\BAR2/BR-7-4/$1I2700/$1N2216 )
  );
  X_BUF   \BAR2/BR-7-4/$1I2700/L  (
    .I(\BAR2/BR-7-4/$1I2700/$1N2216 ),
    .O(\BAR2/BR-7-4/$1N2701 )
  );
  X_ZERO   \BAR2/BR-7-4/$1I2705/$1I2218  (
    .O(\BAR2/BR-7-4/$1I2705/$1N2216 )
  );
  X_BUF   \BAR2/BR-7-4/$1I2705/L  (
    .I(\BAR2/BR-7-4/$1I2705/$1N2216 ),
    .O(\BAR2/BR-7-4/$1N2706 )
  );
  X_OR2   \BAR2/$1I3440/$1I38  (
    .I0(\BAR2/$1I3440/M1 ),
    .I1(\BAR2/$1I3440/M0 ),
    .O(\BAR2/CSREN32 )
  );
  X_AND3   \BAR2/$1I3440/$1I31  (
    .I0(\NlwInverterSignal_BAR2/$1I3440/$1I31/I0 ),
    .I1(CFG74),
    .I2(NlwRenamedSig_OI_CSR1),
    .O(\BAR2/$1I3440/M0 )
  );
  X_AND3   \BAR2/$1I3440/$1I30  (
    .I0(NlwRenamedSig_OI_CSR0),
    .I1(CFG74),
    .I2(CFG110),
    .O(\BAR2/$1I3440/M1 )
  );
  X_OR2   \BAR2/$1I3453/$1I38  (
    .I0(\BAR2/$1I3453/M1 ),
    .I1(\BAR2/$1I3453/M0 ),
    .O(\BAR2/CSREN64 )
  );
  X_AND3   \BAR2/$1I3453/$1I31  (
    .I0(\NlwInverterSignal_BAR2/$1I3453/$1I31/I0 ),
    .I1(CFG74),
    .I2(NlwRenamedSig_OI_CSR1),
    .O(\BAR2/$1I3453/M0 )
  );
  X_AND3   \BAR2/$1I3453/$1I30  (
    .I0(\BAR2/$1N3458 ),
    .I1(CFG74),
    .I2(CFG110),
    .O(\BAR2/$1I3453/M1 )
  );
  X_ZERO   \BAR2/$1I3468/$1I2218  (
    .O(\BAR2/$1I3468/$1N2216 )
  );
  X_BUF   \BAR2/$1I3468/L  (
    .I(\BAR2/$1I3468/$1N2216 ),
    .O(\BAR2/$1N3458 )
  );
  X_ONE   \BAR2/$1I3469/$1I2220  (
    .O(\BAR2/$1I3469/$1N2216 )
  );
  X_BUF   \BAR2/$1I3469/H  (
    .I(\BAR2/$1I3469/$1N2216 ),
    .O(\BAR2/ENABLE32 )
  );
  X_ONE   \BAR2/$2I3304/$1I2220  (
    .O(\BAR2/$2I3304/$1N2216 )
  );
  X_BUF   \BAR2/$2I3304/H  (
    .I(\BAR2/$2I3304/$1N2216 ),
    .O(\BAR2/ENABLENL )
  );
  X_OR2   \BAR2/$2I3321/$1I38  (
    .I0(\BAR2/$2I3321/M1 ),
    .I1(\BAR2/$2I3321/M0 ),
    .O(\BAR2/CSRENNL )
  );
  X_AND3   \BAR2/$2I3321/$1I31  (
    .I0(\NlwInverterSignal_BAR2/$2I3321/$1I31/I0 ),
    .I1(CFG74),
    .I2(NlwRenamedSig_OI_CSR1),
    .O(\BAR2/$2I3321/M0 )
  );
  X_AND3   \BAR2/$2I3321/$1I30  (
    .I0(NlwRenamedSig_OI_CSR0),
    .I1(CFG74),
    .I2(CFG110),
    .O(\BAR2/$2I3321/M1 )
  );
  X_TRI   \F/UPPER/T0  (
    .I(IREG16),
    .O(ADIO16),
    .CTL(\NlwInverterSignal_F/UPPER/T0/T )
  );
  X_TRI   \F/UPPER/T1  (
    .I(IREG17),
    .O(ADIO17),
    .CTL(\NlwInverterSignal_F/UPPER/T1/T )
  );
  X_TRI   \F/UPPER/T2  (
    .I(IREG18),
    .O(ADIO18),
    .CTL(\NlwInverterSignal_F/UPPER/T2/T )
  );
  X_TRI   \F/UPPER/T3  (
    .I(IREG19),
    .O(ADIO19),
    .CTL(\NlwInverterSignal_F/UPPER/T3/T )
  );
  X_TRI   \F/UPPER/T4  (
    .I(IREG20),
    .O(ADIO20),
    .CTL(\NlwInverterSignal_F/UPPER/T4/T )
  );
  X_TRI   \F/UPPER/T5  (
    .I(IREG21),
    .O(ADIO21),
    .CTL(\NlwInverterSignal_F/UPPER/T5/T )
  );
  X_TRI   \F/UPPER/T6  (
    .I(IREG22),
    .O(ADIO22),
    .CTL(\NlwInverterSignal_F/UPPER/T6/T )
  );
  X_TRI   \F/UPPER/T7  (
    .I(IREG23),
    .O(ADIO23),
    .CTL(\NlwInverterSignal_F/UPPER/T7/T )
  );
  X_TRI   \F/UPPER/T8  (
    .I(IREG24),
    .O(ADIO24),
    .CTL(\NlwInverterSignal_F/UPPER/T8/T )
  );
  X_TRI   \F/UPPER/T9  (
    .I(IREG25),
    .O(ADIO25),
    .CTL(\NlwInverterSignal_F/UPPER/T9/T )
  );
  X_TRI   \F/UPPER/T10  (
    .I(IREG26),
    .O(ADIO26),
    .CTL(\NlwInverterSignal_F/UPPER/T10/T )
  );
  X_TRI   \F/UPPER/T11  (
    .I(IREG27),
    .O(ADIO27),
    .CTL(\NlwInverterSignal_F/UPPER/T11/T )
  );
  X_TRI   \F/UPPER/T12  (
    .I(IREG28),
    .O(ADIO28),
    .CTL(\NlwInverterSignal_F/UPPER/T12/T )
  );
  X_TRI   \F/UPPER/T13  (
    .I(IREG29),
    .O(ADIO29),
    .CTL(\NlwInverterSignal_F/UPPER/T13/T )
  );
  X_TRI   \F/UPPER/T14  (
    .I(IREG30),
    .O(ADIO30),
    .CTL(\NlwInverterSignal_F/UPPER/T14/T )
  );
  X_TRI   \F/UPPER/T15  (
    .I(IREG31),
    .O(ADIO31),
    .CTL(\NlwInverterSignal_F/UPPER/T15/T )
  );
  X_TRI   \F/LOWER/T0  (
    .I(IREG0),
    .O(ADIO0),
    .CTL(\NlwInverterSignal_F/LOWER/T0/T )
  );
  X_TRI   \F/LOWER/T1  (
    .I(IREG1),
    .O(ADIO1),
    .CTL(\NlwInverterSignal_F/LOWER/T1/T )
  );
  X_TRI   \F/LOWER/T2  (
    .I(IREG2),
    .O(ADIO2),
    .CTL(\NlwInverterSignal_F/LOWER/T2/T )
  );
  X_TRI   \F/LOWER/T3  (
    .I(IREG3),
    .O(ADIO3),
    .CTL(\NlwInverterSignal_F/LOWER/T3/T )
  );
  X_TRI   \F/LOWER/T4  (
    .I(IREG4),
    .O(ADIO4),
    .CTL(\NlwInverterSignal_F/LOWER/T4/T )
  );
  X_TRI   \F/LOWER/T5  (
    .I(IREG5),
    .O(ADIO5),
    .CTL(\NlwInverterSignal_F/LOWER/T5/T )
  );
  X_TRI   \F/LOWER/T6  (
    .I(IREG6),
    .O(ADIO6),
    .CTL(\NlwInverterSignal_F/LOWER/T6/T )
  );
  X_TRI   \F/LOWER/T7  (
    .I(IREG7),
    .O(ADIO7),
    .CTL(\NlwInverterSignal_F/LOWER/T7/T )
  );
  X_TRI   \F/LOWER/T8  (
    .I(IREG8),
    .O(ADIO8),
    .CTL(\NlwInverterSignal_F/LOWER/T8/T )
  );
  X_TRI   \F/LOWER/T9  (
    .I(IREG9),
    .O(ADIO9),
    .CTL(\NlwInverterSignal_F/LOWER/T9/T )
  );
  X_TRI   \F/LOWER/T10  (
    .I(IREG10),
    .O(ADIO10),
    .CTL(\NlwInverterSignal_F/LOWER/T10/T )
  );
  X_TRI   \F/LOWER/T11  (
    .I(IREG11),
    .O(ADIO11),
    .CTL(\NlwInverterSignal_F/LOWER/T11/T )
  );
  X_TRI   \F/LOWER/T12  (
    .I(IREG12),
    .O(ADIO12),
    .CTL(\NlwInverterSignal_F/LOWER/T12/T )
  );
  X_TRI   \F/LOWER/T13  (
    .I(IREG13),
    .O(ADIO13),
    .CTL(\NlwInverterSignal_F/LOWER/T13/T )
  );
  X_TRI   \F/LOWER/T14  (
    .I(IREG14),
    .O(ADIO14),
    .CTL(\NlwInverterSignal_F/LOWER/T14/T )
  );
  X_TRI   \F/LOWER/T15  (
    .I(IREG15),
    .O(ADIO15),
    .CTL(\NlwInverterSignal_F/LOWER/T15/T )
  );
  X_TRI   \1/UPPER/T0  (
    .I(NlwRenamedSig_OI_CSR16),
    .O(ADIO16),
    .CTL(\NlwInverterSignal_1/UPPER/T0/T )
  );
  X_TRI   \1/UPPER/T1  (
    .I(NlwRenamedSig_OI_CSR17),
    .O(ADIO17),
    .CTL(\NlwInverterSignal_1/UPPER/T1/T )
  );
  X_TRI   \1/UPPER/T2  (
    .I(NlwRenamedSig_OI_CSR18),
    .O(ADIO18),
    .CTL(\NlwInverterSignal_1/UPPER/T2/T )
  );
  X_TRI   \1/UPPER/T3  (
    .I(NlwRenamedSig_OI_CSR19),
    .O(ADIO19),
    .CTL(\NlwInverterSignal_1/UPPER/T3/T )
  );
  X_TRI   \1/UPPER/T4  (
    .I(NlwRenamedSig_OI_CSR20),
    .O(ADIO20),
    .CTL(\NlwInverterSignal_1/UPPER/T4/T )
  );
  X_TRI   \1/UPPER/T5  (
    .I(NlwRenamedSig_OI_CSR21),
    .O(ADIO21),
    .CTL(\NlwInverterSignal_1/UPPER/T5/T )
  );
  X_TRI   \1/UPPER/T6  (
    .I(NlwRenamedSig_OI_CSR22),
    .O(ADIO22),
    .CTL(\NlwInverterSignal_1/UPPER/T6/T )
  );
  X_TRI   \1/UPPER/T7  (
    .I(NlwRenamedSig_OI_CSR23),
    .O(ADIO23),
    .CTL(\NlwInverterSignal_1/UPPER/T7/T )
  );
  X_TRI   \1/UPPER/T8  (
    .I(NlwRenamedSig_OI_CSR24),
    .O(ADIO24),
    .CTL(\NlwInverterSignal_1/UPPER/T8/T )
  );
  X_TRI   \1/UPPER/T9  (
    .I(NlwRenamedSig_OI_CSR25),
    .O(ADIO25),
    .CTL(\NlwInverterSignal_1/UPPER/T9/T )
  );
  X_TRI   \1/UPPER/T10  (
    .I(NlwRenamedSig_OI_CSR26),
    .O(ADIO26),
    .CTL(\NlwInverterSignal_1/UPPER/T10/T )
  );
  X_TRI   \1/UPPER/T11  (
    .I(NlwRenamedSig_OI_CSR27),
    .O(ADIO27),
    .CTL(\NlwInverterSignal_1/UPPER/T11/T )
  );
  X_TRI   \1/UPPER/T12  (
    .I(NlwRenamedSig_OI_CSR28),
    .O(ADIO28),
    .CTL(\NlwInverterSignal_1/UPPER/T12/T )
  );
  X_TRI   \1/UPPER/T13  (
    .I(NlwRenamedSig_OI_CSR29),
    .O(ADIO29),
    .CTL(\NlwInverterSignal_1/UPPER/T13/T )
  );
  X_TRI   \1/UPPER/T14  (
    .I(NlwRenamedSig_OI_CSR30),
    .O(ADIO30),
    .CTL(\NlwInverterSignal_1/UPPER/T14/T )
  );
  X_TRI   \1/UPPER/T15  (
    .I(NlwRenamedSig_OI_CSR31),
    .O(ADIO31),
    .CTL(\NlwInverterSignal_1/UPPER/T15/T )
  );
  X_TRI   \1/LOWER/T0  (
    .I(NlwRenamedSig_OI_CSR0),
    .O(ADIO0),
    .CTL(\NlwInverterSignal_1/LOWER/T0/T )
  );
  X_TRI   \1/LOWER/T1  (
    .I(NlwRenamedSig_OI_CSR1),
    .O(ADIO1),
    .CTL(\NlwInverterSignal_1/LOWER/T1/T )
  );
  X_TRI   \1/LOWER/T2  (
    .I(NlwRenamedSig_OI_CSR2),
    .O(ADIO2),
    .CTL(\NlwInverterSignal_1/LOWER/T2/T )
  );
  X_TRI   \1/LOWER/T3  (
    .I(NlwRenamedSig_OI_CSR3),
    .O(ADIO3),
    .CTL(\NlwInverterSignal_1/LOWER/T3/T )
  );
  X_TRI   \1/LOWER/T4  (
    .I(NlwRenamedSig_OI_CSR4),
    .O(ADIO4),
    .CTL(\NlwInverterSignal_1/LOWER/T4/T )
  );
  X_TRI   \1/LOWER/T5  (
    .I(NlwRenamedSig_OI_CSR5),
    .O(ADIO5),
    .CTL(\NlwInverterSignal_1/LOWER/T5/T )
  );
  X_TRI   \1/LOWER/T6  (
    .I(NlwRenamedSig_OI_CSR6),
    .O(ADIO6),
    .CTL(\NlwInverterSignal_1/LOWER/T6/T )
  );
  X_TRI   \1/LOWER/T7  (
    .I(NlwRenamedSig_OI_CSR7),
    .O(ADIO7),
    .CTL(\NlwInverterSignal_1/LOWER/T7/T )
  );
  X_TRI   \1/LOWER/T8  (
    .I(NlwRenamedSig_OI_CSR8),
    .O(ADIO8),
    .CTL(\NlwInverterSignal_1/LOWER/T8/T )
  );
  X_TRI   \1/LOWER/T9  (
    .I(NlwRenamedSig_OI_CSR9),
    .O(ADIO9),
    .CTL(\NlwInverterSignal_1/LOWER/T9/T )
  );
  X_TRI   \1/LOWER/T10  (
    .I(NlwRenamedSig_OI_CSR10),
    .O(ADIO10),
    .CTL(\NlwInverterSignal_1/LOWER/T10/T )
  );
  X_TRI   \1/LOWER/T11  (
    .I(NlwRenamedSig_OI_CSR11),
    .O(ADIO11),
    .CTL(\NlwInverterSignal_1/LOWER/T11/T )
  );
  X_TRI   \1/LOWER/T12  (
    .I(NlwRenamedSig_OI_CSR12),
    .O(ADIO12),
    .CTL(\NlwInverterSignal_1/LOWER/T12/T )
  );
  X_TRI   \1/LOWER/T13  (
    .I(NlwRenamedSig_OI_CSR13),
    .O(ADIO13),
    .CTL(\NlwInverterSignal_1/LOWER/T13/T )
  );
  X_TRI   \1/LOWER/T14  (
    .I(NlwRenamedSig_OI_CSR14),
    .O(ADIO14),
    .CTL(\NlwInverterSignal_1/LOWER/T14/T )
  );
  X_TRI   \1/LOWER/T15  (
    .I(NlwRenamedSig_OI_CSR15),
    .O(ADIO15),
    .CTL(\NlwInverterSignal_1/LOWER/T15/T )
  );
  X_TRI   \0/UPPER/T0  (
    .I(MD16),
    .O(ADIO16),
    .CTL(\NlwInverterSignal_0/UPPER/T0/T )
  );
  X_TRI   \0/UPPER/T1  (
    .I(MD17),
    .O(ADIO17),
    .CTL(\NlwInverterSignal_0/UPPER/T1/T )
  );
  X_TRI   \0/UPPER/T2  (
    .I(MD18),
    .O(ADIO18),
    .CTL(\NlwInverterSignal_0/UPPER/T2/T )
  );
  X_TRI   \0/UPPER/T3  (
    .I(MD19),
    .O(ADIO19),
    .CTL(\NlwInverterSignal_0/UPPER/T3/T )
  );
  X_TRI   \0/UPPER/T4  (
    .I(MD20),
    .O(ADIO20),
    .CTL(\NlwInverterSignal_0/UPPER/T4/T )
  );
  X_TRI   \0/UPPER/T5  (
    .I(MD21),
    .O(ADIO21),
    .CTL(\NlwInverterSignal_0/UPPER/T5/T )
  );
  X_TRI   \0/UPPER/T6  (
    .I(MD22),
    .O(ADIO22),
    .CTL(\NlwInverterSignal_0/UPPER/T6/T )
  );
  X_TRI   \0/UPPER/T7  (
    .I(MD23),
    .O(ADIO23),
    .CTL(\NlwInverterSignal_0/UPPER/T7/T )
  );
  X_TRI   \0/UPPER/T8  (
    .I(MD24),
    .O(ADIO24),
    .CTL(\NlwInverterSignal_0/UPPER/T8/T )
  );
  X_TRI   \0/UPPER/T9  (
    .I(MD25),
    .O(ADIO25),
    .CTL(\NlwInverterSignal_0/UPPER/T9/T )
  );
  X_TRI   \0/UPPER/T10  (
    .I(MD26),
    .O(ADIO26),
    .CTL(\NlwInverterSignal_0/UPPER/T10/T )
  );
  X_TRI   \0/UPPER/T11  (
    .I(MD27),
    .O(ADIO27),
    .CTL(\NlwInverterSignal_0/UPPER/T11/T )
  );
  X_TRI   \0/UPPER/T12  (
    .I(MD28),
    .O(ADIO28),
    .CTL(\NlwInverterSignal_0/UPPER/T12/T )
  );
  X_TRI   \0/UPPER/T13  (
    .I(MD29),
    .O(ADIO29),
    .CTL(\NlwInverterSignal_0/UPPER/T13/T )
  );
  X_TRI   \0/UPPER/T14  (
    .I(MD30),
    .O(ADIO30),
    .CTL(\NlwInverterSignal_0/UPPER/T14/T )
  );
  X_TRI   \0/UPPER/T15  (
    .I(MD31),
    .O(ADIO31),
    .CTL(\NlwInverterSignal_0/UPPER/T15/T )
  );
  X_TRI   \0/LOWER/T0  (
    .I(MD0),
    .O(ADIO0),
    .CTL(\NlwInverterSignal_0/LOWER/T0/T )
  );
  X_TRI   \0/LOWER/T1  (
    .I(MD1),
    .O(ADIO1),
    .CTL(\NlwInverterSignal_0/LOWER/T1/T )
  );
  X_TRI   \0/LOWER/T2  (
    .I(MD2),
    .O(ADIO2),
    .CTL(\NlwInverterSignal_0/LOWER/T2/T )
  );
  X_TRI   \0/LOWER/T3  (
    .I(MD3),
    .O(ADIO3),
    .CTL(\NlwInverterSignal_0/LOWER/T3/T )
  );
  X_TRI   \0/LOWER/T4  (
    .I(MD4),
    .O(ADIO4),
    .CTL(\NlwInverterSignal_0/LOWER/T4/T )
  );
  X_TRI   \0/LOWER/T5  (
    .I(MD5),
    .O(ADIO5),
    .CTL(\NlwInverterSignal_0/LOWER/T5/T )
  );
  X_TRI   \0/LOWER/T6  (
    .I(MD6),
    .O(ADIO6),
    .CTL(\NlwInverterSignal_0/LOWER/T6/T )
  );
  X_TRI   \0/LOWER/T7  (
    .I(MD7),
    .O(ADIO7),
    .CTL(\NlwInverterSignal_0/LOWER/T7/T )
  );
  X_TRI   \0/LOWER/T8  (
    .I(MD8),
    .O(ADIO8),
    .CTL(\NlwInverterSignal_0/LOWER/T8/T )
  );
  X_TRI   \0/LOWER/T9  (
    .I(MD9),
    .O(ADIO9),
    .CTL(\NlwInverterSignal_0/LOWER/T9/T )
  );
  X_TRI   \0/LOWER/T10  (
    .I(MD10),
    .O(ADIO10),
    .CTL(\NlwInverterSignal_0/LOWER/T10/T )
  );
  X_TRI   \0/LOWER/T11  (
    .I(MD11),
    .O(ADIO11),
    .CTL(\NlwInverterSignal_0/LOWER/T11/T )
  );
  X_TRI   \0/LOWER/T12  (
    .I(MD12),
    .O(ADIO12),
    .CTL(\NlwInverterSignal_0/LOWER/T12/T )
  );
  X_TRI   \0/LOWER/T13  (
    .I(MD13),
    .O(ADIO13),
    .CTL(\NlwInverterSignal_0/LOWER/T13/T )
  );
  X_TRI   \0/LOWER/T14  (
    .I(MD14),
    .O(ADIO14),
    .CTL(\NlwInverterSignal_0/LOWER/T14/T )
  );
  X_TRI   \0/LOWER/T15  (
    .I(MD15),
    .O(ADIO15),
    .CTL(\NlwInverterSignal_0/LOWER/T15/T )
  );
  X_BUF   \PCI-IREG/$1I2604  (
    .I(CFG216),
    .O(IREG16)
  );
  X_BUF   \PCI-IREG/$1I2603  (
    .I(CFG217),
    .O(IREG17)
  );
  X_BUF   \PCI-IREG/$1I2602  (
    .I(CFG218),
    .O(IREG18)
  );
  X_BUF   \PCI-IREG/$1I2601  (
    .I(CFG219),
    .O(IREG19)
  );
  X_BUF   \PCI-IREG/$1I2600  (
    .I(CFG220),
    .O(IREG20)
  );
  X_BUF   \PCI-IREG/$1I2599  (
    .I(CFG221),
    .O(IREG21)
  );
  X_BUF   \PCI-IREG/$1I2598  (
    .I(CFG222),
    .O(IREG22)
  );
  X_BUF   \PCI-IREG/$1I2597  (
    .I(CFG223),
    .O(IREG23)
  );
  X_BUF   \PCI-IREG/$1I2596  (
    .I(CFG224),
    .O(IREG24)
  );
  X_BUF   \PCI-IREG/$1I2595  (
    .I(CFG225),
    .O(IREG25)
  );
  X_BUF   \PCI-IREG/$1I2594  (
    .I(CFG226),
    .O(IREG26)
  );
  X_BUF   \PCI-IREG/$1I2593  (
    .I(CFG227),
    .O(IREG27)
  );
  X_BUF   \PCI-IREG/$1I2592  (
    .I(CFG228),
    .O(IREG28)
  );
  X_BUF   \PCI-IREG/$1I2591  (
    .I(CFG229),
    .O(IREG29)
  );
  X_BUF   \PCI-IREG/$1I2590  (
    .I(CFG230),
    .O(IREG30)
  );
  X_BUF   \PCI-IREG/$1I2589  (
    .I(CFG231),
    .O(IREG31)
  );
  X_BUF   \PCI-IREG/INT-PINX/$1I2499  (
    .I(CFG113),
    .O(IREG8)
  );
  X_ZERO   \PCI-IREG/INT-PINX/$1I2486/$1I2218  (
    .O(\PCI-IREG/INT-PINX/$1I2486/$1N2216 )
  );
  X_BUF   \PCI-IREG/INT-PINX/$1I2486/L  (
    .I(\PCI-IREG/INT-PINX/$1I2486/$1N2216 ),
    .O(IREG9)
  );
  X_ZERO   \PCI-IREG/INT-PINX/$1I2488/$1I2218  (
    .O(\PCI-IREG/INT-PINX/$1I2488/$1N2216 )
  );
  X_BUF   \PCI-IREG/INT-PINX/$1I2488/L  (
    .I(\PCI-IREG/INT-PINX/$1I2488/$1N2216 ),
    .O(IREG10)
  );
  X_ZERO   \PCI-IREG/INT-PINX/$1I2490/$1I2218  (
    .O(\PCI-IREG/INT-PINX/$1I2490/$1N2216 )
  );
  X_BUF   \PCI-IREG/INT-PINX/$1I2490/L  (
    .I(\PCI-IREG/INT-PINX/$1I2490/$1N2216 ),
    .O(IREG11)
  );
  X_ZERO   \PCI-IREG/INT-PINX/$1I2492/$1I2218  (
    .O(\PCI-IREG/INT-PINX/$1I2492/$1N2216 )
  );
  X_BUF   \PCI-IREG/INT-PINX/$1I2492/L  (
    .I(\PCI-IREG/INT-PINX/$1I2492/$1N2216 ),
    .O(IREG12)
  );
  X_ZERO   \PCI-IREG/INT-PINX/$1I2494/$1I2218  (
    .O(\PCI-IREG/INT-PINX/$1I2494/$1N2216 )
  );
  X_BUF   \PCI-IREG/INT-PINX/$1I2494/L  (
    .I(\PCI-IREG/INT-PINX/$1I2494/$1N2216 ),
    .O(IREG13)
  );
  X_ZERO   \PCI-IREG/INT-PINX/$1I2496/$1I2218  (
    .O(\PCI-IREG/INT-PINX/$1I2496/$1N2216 )
  );
  X_BUF   \PCI-IREG/INT-PINX/$1I2496/L  (
    .I(\PCI-IREG/INT-PINX/$1I2496/$1N2216 ),
    .O(IREG14)
  );
  X_ZERO   \PCI-IREG/INT-PINX/$1I2498/$1I2218  (
    .O(\PCI-IREG/INT-PINX/$1I2498/$1N2216 )
  );
  X_BUF   \PCI-IREG/INT-PINX/$1I2498/L  (
    .I(\PCI-IREG/INT-PINX/$1I2498/$1N2216 ),
    .O(IREG15)
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-IREG/INT-LNX/Q7  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(CE15_0),
    .CLK(CLK),
    .I(ADIO7),
    .O(IREG7),
    .RST(GND)
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-IREG/INT-LNX/Q1  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(CE15_0),
    .CLK(CLK),
    .I(ADIO1),
    .O(IREG1),
    .RST(GND)
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-IREG/INT-LNX/Q5  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(CE15_0),
    .CLK(CLK),
    .I(ADIO5),
    .O(IREG5),
    .RST(GND)
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-IREG/INT-LNX/Q3  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(CE15_0),
    .CLK(CLK),
    .I(ADIO3),
    .O(IREG3),
    .RST(GND)
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-IREG/INT-LNX/Q0  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(CE15_0),
    .CLK(CLK),
    .I(ADIO0),
    .O(IREG0),
    .RST(GND)
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-IREG/INT-LNX/Q2  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(CE15_0),
    .CLK(CLK),
    .I(ADIO2),
    .O(IREG2),
    .RST(GND)
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-IREG/INT-LNX/Q4  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(CE15_0),
    .CLK(CLK),
    .I(ADIO4),
    .O(IREG4),
    .RST(GND)
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-IREG/INT-LNX/Q6  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(CE15_0),
    .CLK(CLK),
    .I(ADIO6),
    .O(IREG6),
    .RST(GND)
  );
  X_BUF   \PCI-IREG/$1I2521/NC  (
    .I(CE15_1),
    .O(\NLW_PCI-IREG/$1I2521/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-IREG/$1I2555/NC  (
    .I(ADIO15),
    .O(\NLW_PCI-IREG/$1I2555/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-IREG/$1I2557/NC  (
    .I(ADIO14),
    .O(\NLW_PCI-IREG/$1I2557/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-IREG/$1I2559/NC  (
    .I(ADIO13),
    .O(\NLW_PCI-IREG/$1I2559/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-IREG/$1I2561/NC  (
    .I(ADIO12),
    .O(\NLW_PCI-IREG/$1I2561/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-IREG/$1I2563/NC  (
    .I(ADIO11),
    .O(\NLW_PCI-IREG/$1I2563/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-IREG/$1I2565/NC  (
    .I(ADIO10),
    .O(\NLW_PCI-IREG/$1I2565/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-IREG/$1I2567/NC  (
    .I(ADIO9),
    .O(\NLW_PCI-IREG/$1I2567/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-IREG/$1I2569/NC  (
    .I(ADIO8),
    .O(\NLW_PCI-IREG/$1I2569/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-IREG/$1I2582/NC  (
    .I(CE15_2),
    .O(\NLW_PCI-IREG/$1I2582/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-IREG/$1I2584/NC  (
    .I(CE15_3),
    .O(\NLW_PCI-IREG/$1I2584/NC_O_UNCONNECTED )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CSR/CMDREG/Q10  (
    .CE(CE1_1),
    .CLK(CLK),
    .I(ADIO10),
    .O(NlwRenamedSig_OI_CSR10),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND2   \PCI-CSR/CMDREG/$1I2564  (
    .I0(HAS_IO),
    .I1(\PCI-CSR/CMDREG/$1N2346 ),
    .O(NlwRenamedSig_OI_CSR0)
  );
  X_AND2   \PCI-CSR/CMDREG/$1I2563  (
    .I0(HAS_MEM),
    .I1(\PCI-CSR/CMDREG/$1N2446 ),
    .O(NlwRenamedSig_OI_CSR1)
  );
  X_BUF   \PCI-CSR/CMDREG/$1I2535  (
    .I(\PCI-CSR/CMDREG/$1N2560 ),
    .O(NlwRenamedSig_OI_CSR5)
  );
  X_BUF   \PCI-CSR/CMDREG/$1I2511  (
    .I(\PCI-CSR/CMDREG/$1N2556 ),
    .O(NlwRenamedSig_OI_CSR3)
  );
  X_BUF   \PCI-CSR/CMDREG/$1I2488  (
    .I(\PCI-CSR/CMDREG/$1N2562 ),
    .O(NlwRenamedSig_OI_CSR7)
  );
  X_BUF   \PCI-CSR/CMDREG/$1I2483  (
    .I(\PCI-CSR/CMDREG/$1N2559 ),
    .O(NlwRenamedSig_OI_CSR4)
  );
  X_BUF   \PCI-CSR/CMDREG/$1I2479  (
    .I(\PCI-CSR/CMDREG/$1N2514 ),
    .O(NlwRenamedSig_OI_CSR15)
  );
  X_BUF   \PCI-CSR/CMDREG/$1I2471  (
    .I(\PCI-CSR/CMDREG/$1N2527 ),
    .O(NlwRenamedSig_OI_CSR9)
  );
  X_BUF   \PCI-CSR/CMDREG/$1I2470  (
    .I(\PCI-CSR/CMDREG/$1N2524 ),
    .O(NlwRenamedSig_OI_CSR11)
  );
  X_BUF   \PCI-CSR/CMDREG/$1I2469  (
    .I(\PCI-CSR/CMDREG/$1N2525 ),
    .O(NlwRenamedSig_OI_CSR12)
  );
  X_BUF   \PCI-CSR/CMDREG/$1I2468  (
    .I(\PCI-CSR/CMDREG/$1N2523 ),
    .O(NlwRenamedSig_OI_CSR13)
  );
  X_BUF   \PCI-CSR/CMDREG/$1I2467  (
    .I(\PCI-CSR/CMDREG/$1N2522 ),
    .O(NlwRenamedSig_OI_CSR14)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CSR/CMDREG/Q1  (
    .CE(CE1_0),
    .CLK(CLK),
    .I(ADIO1),
    .O(\PCI-CSR/CMDREG/$1N2446 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CSR/CMDREG/Q0  (
    .CE(CE1_0),
    .CLK(CLK),
    .I(ADIO0),
    .O(\PCI-CSR/CMDREG/$1N2346 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CSR/CMDREG/Q8  (
    .CE(CE1_1),
    .CLK(CLK),
    .I(ADIO8),
    .O(NlwRenamedSig_OI_CSR8),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CSR/CMDREG/Q2  (
    .CE(CE1_0),
    .CLK(CLK),
    .I(ADIO2),
    .O(NlwRenamedSig_OI_CSR2),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CSR/CMDREG/Q6  (
    .CE(CE1_0),
    .CLK(CLK),
    .I(ADIO6),
    .O(NlwRenamedSig_OI_CSR6),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_BUF   \PCI-CSR/CMDREG/$1I2492/NC  (
    .I(ADIO15),
    .O(\NLW_PCI-CSR/CMDREG/$1I2492/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-CSR/CMDREG/$1I2495/NC  (
    .I(ADIO14),
    .O(\NLW_PCI-CSR/CMDREG/$1I2495/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-CSR/CMDREG/$1I2497/NC  (
    .I(ADIO13),
    .O(\NLW_PCI-CSR/CMDREG/$1I2497/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-CSR/CMDREG/$1I2499/NC  (
    .I(ADIO12),
    .O(\NLW_PCI-CSR/CMDREG/$1I2499/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-CSR/CMDREG/$1I2501/NC  (
    .I(ADIO11),
    .O(\NLW_PCI-CSR/CMDREG/$1I2501/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-CSR/CMDREG/$1I2505/NC  (
    .I(ADIO9),
    .O(\NLW_PCI-CSR/CMDREG/$1I2505/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-CSR/CMDREG/$1I2507/NC  (
    .I(ADIO7),
    .O(\NLW_PCI-CSR/CMDREG/$1I2507/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-CSR/CMDREG/$1I2509/NC  (
    .I(ADIO5),
    .O(\NLW_PCI-CSR/CMDREG/$1I2509/NC_O_UNCONNECTED )
  );
  X_ZERO   \PCI-CSR/CMDREG/$1I2520/$1I2218  (
    .O(\PCI-CSR/CMDREG/$1I2520/$1N2216 )
  );
  X_BUF   \PCI-CSR/CMDREG/$1I2520/L  (
    .I(\PCI-CSR/CMDREG/$1I2520/$1N2216 ),
    .O(\PCI-CSR/CMDREG/$1N2514 )
  );
  X_ZERO   \PCI-CSR/CMDREG/$1I2521/$1I2218  (
    .O(\PCI-CSR/CMDREG/$1I2521/$1N2216 )
  );
  X_BUF   \PCI-CSR/CMDREG/$1I2521/L  (
    .I(\PCI-CSR/CMDREG/$1I2521/$1N2216 ),
    .O(\PCI-CSR/CMDREG/$1N2522 )
  );
  X_ZERO   \PCI-CSR/CMDREG/$1I2528/$1I2218  (
    .O(\PCI-CSR/CMDREG/$1I2528/$1N2216 )
  );
  X_BUF   \PCI-CSR/CMDREG/$1I2528/L  (
    .I(\PCI-CSR/CMDREG/$1I2528/$1N2216 ),
    .O(\PCI-CSR/CMDREG/$1N2523 )
  );
  X_ZERO   \PCI-CSR/CMDREG/$1I2529/$1I2218  (
    .O(\PCI-CSR/CMDREG/$1I2529/$1N2216 )
  );
  X_BUF   \PCI-CSR/CMDREG/$1I2529/L  (
    .I(\PCI-CSR/CMDREG/$1I2529/$1N2216 ),
    .O(\PCI-CSR/CMDREG/$1N2525 )
  );
  X_ZERO   \PCI-CSR/CMDREG/$1I2530/$1I2218  (
    .O(\PCI-CSR/CMDREG/$1I2530/$1N2216 )
  );
  X_BUF   \PCI-CSR/CMDREG/$1I2530/L  (
    .I(\PCI-CSR/CMDREG/$1I2530/$1N2216 ),
    .O(\PCI-CSR/CMDREG/$1N2524 )
  );
  X_ZERO   \PCI-CSR/CMDREG/$1I2532/$1I2218  (
    .O(\PCI-CSR/CMDREG/$1I2532/$1N2216 )
  );
  X_BUF   \PCI-CSR/CMDREG/$1I2532/L  (
    .I(\PCI-CSR/CMDREG/$1I2532/$1N2216 ),
    .O(\PCI-CSR/CMDREG/$1N2527 )
  );
  X_BUF   \PCI-CSR/CMDREG/$1I2538/NC  (
    .I(ADIO4),
    .O(\NLW_PCI-CSR/CMDREG/$1I2538/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-CSR/CMDREG/$1I2540/NC  (
    .I(ADIO3),
    .O(\NLW_PCI-CSR/CMDREG/$1I2540/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-CSR/CMDREG/$1I2551/NC  (
    .I(CE1_1),
    .O(\NLW_PCI-CSR/CMDREG/$1I2551/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-CSR/CMDREG/$1I2552/NC  (
    .I(CE1_0),
    .O(\NLW_PCI-CSR/CMDREG/$1I2552/NC_O_UNCONNECTED )
  );
  X_ZERO   \PCI-CSR/CMDREG/$1I2557/$1I2218  (
    .O(\PCI-CSR/CMDREG/$1I2557/$1N2216 )
  );
  X_BUF   \PCI-CSR/CMDREG/$1I2557/L  (
    .I(\PCI-CSR/CMDREG/$1I2557/$1N2216 ),
    .O(\PCI-CSR/CMDREG/$1N2556 )
  );
  X_ZERO   \PCI-CSR/CMDREG/$1I2558/$1I2218  (
    .O(\PCI-CSR/CMDREG/$1I2558/$1N2216 )
  );
  X_BUF   \PCI-CSR/CMDREG/$1I2558/L  (
    .I(\PCI-CSR/CMDREG/$1I2558/$1N2216 ),
    .O(\PCI-CSR/CMDREG/$1N2559 )
  );
  X_ZERO   \PCI-CSR/CMDREG/$1I2561/$1I2218  (
    .O(\PCI-CSR/CMDREG/$1I2561/$1N2216 )
  );
  X_BUF   \PCI-CSR/CMDREG/$1I2561/L  (
    .I(\PCI-CSR/CMDREG/$1I2561/$1N2216 ),
    .O(\PCI-CSR/CMDREG/$1N2560 )
  );
  X_ZERO   \PCI-CSR/CMDREG/$1I2583/$1I2218  (
    .O(\PCI-CSR/CMDREG/$1I2583/$1N2216 )
  );
  X_BUF   \PCI-CSR/CMDREG/$1I2583/L  (
    .I(\PCI-CSR/CMDREG/$1I2583/$1N2216 ),
    .O(\PCI-CSR/CMDREG/$1N2562 )
  );
  X_INV   \PCI-CSR/STATREG/$1I2632  (
    .I(INTR_N),
    .O(\PCI-CSR/STATREG/$1N2634 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CSR/STATREG/$1I2627  (
    .CE(\PCI-CSR/STATREG/$1N2630 ),
    .CLK(CLK),
    .I(\PCI-CSR/STATREG/$1N2634 ),
    .O(NlwRenamedSig_OI_CSR19),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_BUF   \PCI-CSR/STATREG/$1I2593  (
    .I(\PCI-CSR/STATREG/$1N2595 ),
    .O(NlwRenamedSig_OI_CSR22)
  );
  X_BUF   \PCI-CSR/STATREG/$1I2589  (
    .I(\PCI-CSR/STATREG/$1N2588 ),
    .O(NlwRenamedSig_OI_CSR25)
  );
  X_BUF   \PCI-CSR/STATREG/$1I2586  (
    .I(\PCI-CSR/STATREG/$1N2585 ),
    .O(NlwRenamedSig_OI_CSR26)
  );
  X_BUF   \PCI-CSR/STATREG/$1I2485  (
    .I(\PCI-CSR/STATREG/$1N2474 ),
    .O(NlwRenamedSig_OI_CSR23)
  );
  X_BUF   \PCI-CSR/STATREG/$1I2481  (
    .I(CFG244),
    .O(NlwRenamedSig_OI_CSR21)
  );
  X_BUF   \PCI-CSR/STATREG/$1I2473  (
    .I(CFG116),
    .O(NlwRenamedSig_OI_CSR20)
  );
  X_BUF   \PCI-CSR/STATREG/$1I2471  (
    .I(\PCI-CSR/STATREG/$1N2605 ),
    .O(NlwRenamedSig_OI_CSR18)
  );
  X_BUF   \PCI-CSR/STATREG/$1I2470  (
    .I(\PCI-CSR/STATREG/$1N2606 ),
    .O(NlwRenamedSig_OI_CSR17)
  );
  X_BUF   \PCI-CSR/STATREG/$1I2469  (
    .I(\PCI-CSR/STATREG/$1N2609 ),
    .O(NlwRenamedSig_OI_CSR16)
  );
  X_OR2   \PCI-CSR/STATREG/Q14/$1I2236  (
    .I0(SET14),
    .I1(\PCI-CSR/STATREG/Q14/$1N2238 ),
    .O(\PCI-CSR/STATREG/Q14/D )
  );
  X_AND2   \PCI-CSR/STATREG/Q14/$1I2230  (
    .I0(\NlwInverterSignal_PCI-CSR/STATREG/Q14/$1I2230/I0 ),
    .I1(NlwRenamedSig_OI_CSR30),
    .O(\PCI-CSR/STATREG/Q14/$1N2240 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CSR/STATREG/Q14/FDCE  (
    .CE(VCC),
    .CLK(CLK),
    .I(\PCI-CSR/STATREG/Q14/D ),
    .O(NlwRenamedSig_OI_CSR30),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND2   \PCI-CSR/STATREG/Q14/$1I2233/$1I9  (
    .I0(\PCI-CSR/STATREG/Q14/$1N2240 ),
    .I1(CE1_3),
    .O(\PCI-CSR/STATREG/Q14/$1I2233/M1 )
  );
  X_OR2   \PCI-CSR/STATREG/Q14/$1I2233/$1I8  (
    .I0(\PCI-CSR/STATREG/Q14/$1I2233/M1 ),
    .I1(\PCI-CSR/STATREG/Q14/$1I2233/M0 ),
    .O(\PCI-CSR/STATREG/Q14/$1N2238 )
  );
  X_AND2   \PCI-CSR/STATREG/Q14/$1I2233/$1I7  (
    .I0(\NlwInverterSignal_PCI-CSR/STATREG/Q14/$1I2233/$1I7/I0 ),
    .I1(NlwRenamedSig_OI_CSR30),
    .O(\PCI-CSR/STATREG/Q14/$1I2233/M0 )
  );
  X_OR2   \PCI-CSR/STATREG/Q12/$1I2236  (
    .I0(SET12),
    .I1(\PCI-CSR/STATREG/Q12/$1N2238 ),
    .O(\PCI-CSR/STATREG/Q12/D )
  );
  X_AND2   \PCI-CSR/STATREG/Q12/$1I2230  (
    .I0(\NlwInverterSignal_PCI-CSR/STATREG/Q12/$1I2230/I0 ),
    .I1(NlwRenamedSig_OI_CSR28),
    .O(\PCI-CSR/STATREG/Q12/$1N2240 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CSR/STATREG/Q12/FDCE  (
    .CE(VCC),
    .CLK(CLK),
    .I(\PCI-CSR/STATREG/Q12/D ),
    .O(NlwRenamedSig_OI_CSR28),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND2   \PCI-CSR/STATREG/Q12/$1I2233/$1I9  (
    .I0(\PCI-CSR/STATREG/Q12/$1N2240 ),
    .I1(CE1_3),
    .O(\PCI-CSR/STATREG/Q12/$1I2233/M1 )
  );
  X_OR2   \PCI-CSR/STATREG/Q12/$1I2233/$1I8  (
    .I0(\PCI-CSR/STATREG/Q12/$1I2233/M1 ),
    .I1(\PCI-CSR/STATREG/Q12/$1I2233/M0 ),
    .O(\PCI-CSR/STATREG/Q12/$1N2238 )
  );
  X_AND2   \PCI-CSR/STATREG/Q12/$1I2233/$1I7  (
    .I0(\NlwInverterSignal_PCI-CSR/STATREG/Q12/$1I2233/$1I7/I0 ),
    .I1(NlwRenamedSig_OI_CSR28),
    .O(\PCI-CSR/STATREG/Q12/$1I2233/M0 )
  );
  X_OR2   \PCI-CSR/STATREG/Q8/$1I2236  (
    .I0(SET8),
    .I1(\PCI-CSR/STATREG/Q8/$1N2238 ),
    .O(\PCI-CSR/STATREG/Q8/D )
  );
  X_AND2   \PCI-CSR/STATREG/Q8/$1I2230  (
    .I0(\NlwInverterSignal_PCI-CSR/STATREG/Q8/$1I2230/I0 ),
    .I1(NlwRenamedSig_OI_CSR24),
    .O(\PCI-CSR/STATREG/Q8/$1N2240 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CSR/STATREG/Q8/FDCE  (
    .CE(VCC),
    .CLK(CLK),
    .I(\PCI-CSR/STATREG/Q8/D ),
    .O(NlwRenamedSig_OI_CSR24),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND2   \PCI-CSR/STATREG/Q8/$1I2233/$1I9  (
    .I0(\PCI-CSR/STATREG/Q8/$1N2240 ),
    .I1(CE1_3),
    .O(\PCI-CSR/STATREG/Q8/$1I2233/M1 )
  );
  X_OR2   \PCI-CSR/STATREG/Q8/$1I2233/$1I8  (
    .I0(\PCI-CSR/STATREG/Q8/$1I2233/M1 ),
    .I1(\PCI-CSR/STATREG/Q8/$1I2233/M0 ),
    .O(\PCI-CSR/STATREG/Q8/$1N2238 )
  );
  X_AND2   \PCI-CSR/STATREG/Q8/$1I2233/$1I7  (
    .I0(\NlwInverterSignal_PCI-CSR/STATREG/Q8/$1I2233/$1I7/I0 ),
    .I1(NlwRenamedSig_OI_CSR24),
    .O(\PCI-CSR/STATREG/Q8/$1I2233/M0 )
  );
  X_OR2   \PCI-CSR/STATREG/Q11/$1I2236  (
    .I0(SET11),
    .I1(\PCI-CSR/STATREG/Q11/$1N2238 ),
    .O(\PCI-CSR/STATREG/Q11/D )
  );
  X_AND2   \PCI-CSR/STATREG/Q11/$1I2230  (
    .I0(\NlwInverterSignal_PCI-CSR/STATREG/Q11/$1I2230/I0 ),
    .I1(NlwRenamedSig_OI_CSR27),
    .O(\PCI-CSR/STATREG/Q11/$1N2240 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CSR/STATREG/Q11/FDCE  (
    .CE(VCC),
    .CLK(CLK),
    .I(\PCI-CSR/STATREG/Q11/D ),
    .O(NlwRenamedSig_OI_CSR27),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND2   \PCI-CSR/STATREG/Q11/$1I2233/$1I9  (
    .I0(\PCI-CSR/STATREG/Q11/$1N2240 ),
    .I1(CE1_3),
    .O(\PCI-CSR/STATREG/Q11/$1I2233/M1 )
  );
  X_OR2   \PCI-CSR/STATREG/Q11/$1I2233/$1I8  (
    .I0(\PCI-CSR/STATREG/Q11/$1I2233/M1 ),
    .I1(\PCI-CSR/STATREG/Q11/$1I2233/M0 ),
    .O(\PCI-CSR/STATREG/Q11/$1N2238 )
  );
  X_AND2   \PCI-CSR/STATREG/Q11/$1I2233/$1I7  (
    .I0(\NlwInverterSignal_PCI-CSR/STATREG/Q11/$1I2233/$1I7/I0 ),
    .I1(NlwRenamedSig_OI_CSR27),
    .O(\PCI-CSR/STATREG/Q11/$1I2233/M0 )
  );
  X_OR2   \PCI-CSR/STATREG/Q13/$1I2236  (
    .I0(SET13),
    .I1(\PCI-CSR/STATREG/Q13/$1N2238 ),
    .O(\PCI-CSR/STATREG/Q13/D )
  );
  X_AND2   \PCI-CSR/STATREG/Q13/$1I2230  (
    .I0(\NlwInverterSignal_PCI-CSR/STATREG/Q13/$1I2230/I0 ),
    .I1(NlwRenamedSig_OI_CSR29),
    .O(\PCI-CSR/STATREG/Q13/$1N2240 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CSR/STATREG/Q13/FDCE  (
    .CE(VCC),
    .CLK(CLK),
    .I(\PCI-CSR/STATREG/Q13/D ),
    .O(NlwRenamedSig_OI_CSR29),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND2   \PCI-CSR/STATREG/Q13/$1I2233/$1I9  (
    .I0(\PCI-CSR/STATREG/Q13/$1N2240 ),
    .I1(CE1_3),
    .O(\PCI-CSR/STATREG/Q13/$1I2233/M1 )
  );
  X_OR2   \PCI-CSR/STATREG/Q13/$1I2233/$1I8  (
    .I0(\PCI-CSR/STATREG/Q13/$1I2233/M1 ),
    .I1(\PCI-CSR/STATREG/Q13/$1I2233/M0 ),
    .O(\PCI-CSR/STATREG/Q13/$1N2238 )
  );
  X_AND2   \PCI-CSR/STATREG/Q13/$1I2233/$1I7  (
    .I0(\NlwInverterSignal_PCI-CSR/STATREG/Q13/$1I2233/$1I7/I0 ),
    .I1(NlwRenamedSig_OI_CSR29),
    .O(\PCI-CSR/STATREG/Q13/$1I2233/M0 )
  );
  X_OR2   \PCI-CSR/STATREG/Q15/$1I2236  (
    .I0(SET15),
    .I1(\PCI-CSR/STATREG/Q15/$1N2238 ),
    .O(\PCI-CSR/STATREG/Q15/D )
  );
  X_AND2   \PCI-CSR/STATREG/Q15/$1I2230  (
    .I0(\NlwInverterSignal_PCI-CSR/STATREG/Q15/$1I2230/I0 ),
    .I1(NlwRenamedSig_OI_CSR31),
    .O(\PCI-CSR/STATREG/Q15/$1N2240 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \PCI-CSR/STATREG/Q15/FDCE  (
    .CE(VCC),
    .CLK(CLK),
    .I(\PCI-CSR/STATREG/Q15/D ),
    .O(NlwRenamedSig_OI_CSR31),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND2   \PCI-CSR/STATREG/Q15/$1I2233/$1I9  (
    .I0(\PCI-CSR/STATREG/Q15/$1N2240 ),
    .I1(CE1_3),
    .O(\PCI-CSR/STATREG/Q15/$1I2233/M1 )
  );
  X_OR2   \PCI-CSR/STATREG/Q15/$1I2233/$1I8  (
    .I0(\PCI-CSR/STATREG/Q15/$1I2233/M1 ),
    .I1(\PCI-CSR/STATREG/Q15/$1I2233/M0 ),
    .O(\PCI-CSR/STATREG/Q15/$1N2238 )
  );
  X_AND2   \PCI-CSR/STATREG/Q15/$1I2233/$1I7  (
    .I0(\NlwInverterSignal_PCI-CSR/STATREG/Q15/$1I2233/$1I7/I0 ),
    .I1(NlwRenamedSig_OI_CSR31),
    .O(\PCI-CSR/STATREG/Q15/$1I2233/M0 )
  );
  X_BUF   \PCI-CSR/STATREG/$1I2497/NC  (
    .I(ADIO26),
    .O(\NLW_PCI-CSR/STATREG/$1I2497/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-CSR/STATREG/$1I2500/NC  (
    .I(ADIO25),
    .O(\NLW_PCI-CSR/STATREG/$1I2500/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-CSR/STATREG/$1I2502/NC  (
    .I(ADIO23),
    .O(\NLW_PCI-CSR/STATREG/$1I2502/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-CSR/STATREG/$1I2504/NC  (
    .I(ADIO21),
    .O(\NLW_PCI-CSR/STATREG/$1I2504/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-CSR/STATREG/$1I2506/NC  (
    .I(ADIO20),
    .O(\NLW_PCI-CSR/STATREG/$1I2506/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-CSR/STATREG/$1I2508/NC  (
    .I(ADIO19),
    .O(\NLW_PCI-CSR/STATREG/$1I2508/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-CSR/STATREG/$1I2510/NC  (
    .I(ADIO18),
    .O(\NLW_PCI-CSR/STATREG/$1I2510/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-CSR/STATREG/$1I2512/NC  (
    .I(ADIO17),
    .O(\NLW_PCI-CSR/STATREG/$1I2512/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-CSR/STATREG/$1I2514/NC  (
    .I(ADIO16),
    .O(\NLW_PCI-CSR/STATREG/$1I2514/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-CSR/STATREG/$1I2523/NC  (
    .I(SET10),
    .O(\NLW_PCI-CSR/STATREG/$1I2523/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-CSR/STATREG/$1I2524/NC  (
    .I(SET9),
    .O(\NLW_PCI-CSR/STATREG/$1I2524/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-CSR/STATREG/$1I2525/NC  (
    .I(SET7),
    .O(\NLW_PCI-CSR/STATREG/$1I2525/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-CSR/STATREG/$1I2526/NC  (
    .I(SET5),
    .O(\NLW_PCI-CSR/STATREG/$1I2526/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-CSR/STATREG/$1I2527/NC  (
    .I(SET4),
    .O(\NLW_PCI-CSR/STATREG/$1I2527/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-CSR/STATREG/$1I2528/NC  (
    .I(SET3),
    .O(\NLW_PCI-CSR/STATREG/$1I2528/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-CSR/STATREG/$1I2529/NC  (
    .I(SET2),
    .O(\NLW_PCI-CSR/STATREG/$1I2529/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-CSR/STATREG/$1I2530/NC  (
    .I(SET1),
    .O(\NLW_PCI-CSR/STATREG/$1I2530/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-CSR/STATREG/$1I2532/NC  (
    .I(SET0),
    .O(\NLW_PCI-CSR/STATREG/$1I2532/NC_O_UNCONNECTED )
  );
  X_ZERO   \PCI-CSR/STATREG/$1I2569/$1I2218  (
    .O(\PCI-CSR/STATREG/$1I2569/$1N2216 )
  );
  X_BUF   \PCI-CSR/STATREG/$1I2569/L  (
    .I(\PCI-CSR/STATREG/$1I2569/$1N2216 ),
    .O(\PCI-CSR/STATREG/$1N2474 )
  );
  X_ZERO   \PCI-CSR/STATREG/$1I2587/$1I2218  (
    .O(\PCI-CSR/STATREG/$1I2587/$1N2216 )
  );
  X_BUF   \PCI-CSR/STATREG/$1I2587/L  (
    .I(\PCI-CSR/STATREG/$1I2587/$1N2216 ),
    .O(\PCI-CSR/STATREG/$1N2585 )
  );
  X_ONE   \PCI-CSR/STATREG/$1I2590/$1I2220  (
    .O(\PCI-CSR/STATREG/$1I2590/$1N2216 )
  );
  X_BUF   \PCI-CSR/STATREG/$1I2590/H  (
    .I(\PCI-CSR/STATREG/$1I2590/$1N2216 ),
    .O(\PCI-CSR/STATREG/$1N2588 )
  );
  X_ZERO   \PCI-CSR/STATREG/$1I2596/$1I2218  (
    .O(\PCI-CSR/STATREG/$1I2596/$1N2216 )
  );
  X_BUF   \PCI-CSR/STATREG/$1I2596/L  (
    .I(\PCI-CSR/STATREG/$1I2596/$1N2216 ),
    .O(\PCI-CSR/STATREG/$1N2595 )
  );
  X_BUF   \PCI-CSR/STATREG/$1I2598/NC  (
    .I(SET6),
    .O(\NLW_PCI-CSR/STATREG/$1I2598/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-CSR/STATREG/$1I2600/NC  (
    .I(ADIO22),
    .O(\NLW_PCI-CSR/STATREG/$1I2600/NC_O_UNCONNECTED )
  );
  X_ZERO   \PCI-CSR/STATREG/$1I2604/$1I2218  (
    .O(\PCI-CSR/STATREG/$1I2604/$1N2216 )
  );
  X_BUF   \PCI-CSR/STATREG/$1I2604/L  (
    .I(\PCI-CSR/STATREG/$1I2604/$1N2216 ),
    .O(\PCI-CSR/STATREG/$1N2605 )
  );
  X_ZERO   \PCI-CSR/STATREG/$1I2607/$1I2218  (
    .O(\PCI-CSR/STATREG/$1I2607/$1N2216 )
  );
  X_BUF   \PCI-CSR/STATREG/$1I2607/L  (
    .I(\PCI-CSR/STATREG/$1I2607/$1N2216 ),
    .O(\PCI-CSR/STATREG/$1N2606 )
  );
  X_ZERO   \PCI-CSR/STATREG/$1I2608/$1I2218  (
    .O(\PCI-CSR/STATREG/$1I2608/$1N2216 )
  );
  X_BUF   \PCI-CSR/STATREG/$1I2608/L  (
    .I(\PCI-CSR/STATREG/$1I2608/$1N2216 ),
    .O(\PCI-CSR/STATREG/$1N2609 )
  );
  X_BUF   \PCI-CSR/STATREG/$1I2612/NC  (
    .I(CE1_3),
    .O(\NLW_PCI-CSR/STATREG/$1I2612/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-CSR/STATREG/$1I2613/NC  (
    .I(CE1_2),
    .O(\NLW_PCI-CSR/STATREG/$1I2613/NC_O_UNCONNECTED )
  );
  X_ONE   \PCI-CSR/STATREG/$1I2631/$1I2220  (
    .O(\PCI-CSR/STATREG/$1I2631/$1N2216 )
  );
  X_BUF   \PCI-CSR/STATREG/$1I2631/H  (
    .I(\PCI-CSR/STATREG/$1I2631/$1N2216 ),
    .O(\PCI-CSR/STATREG/$1N2630 )
  );
  X_OR4   \PCI-ROM/$1I8593  (
    .I0(\PCI-ROM/RA0 ),
    .I1(\PCI-ROM/RB0 ),
    .I2(\PCI-ROM/RE0 ),
    .I3(\PCI-ROM/ROM0 ),
    .O(MD0)
  );
  X_OR4   \PCI-ROM/$1I8592  (
    .I0(\PCI-ROM/RA1 ),
    .I1(\PCI-ROM/RB1 ),
    .I2(\PCI-ROM/RE1 ),
    .I3(\PCI-ROM/ROM1 ),
    .O(MD1)
  );
  X_OR4   \PCI-ROM/$1I8591  (
    .I0(\PCI-ROM/RA2 ),
    .I1(\PCI-ROM/RB2 ),
    .I2(\PCI-ROM/RE2 ),
    .I3(\PCI-ROM/ROM2 ),
    .O(MD2)
  );
  X_OR4   \PCI-ROM/$1I8590  (
    .I0(\PCI-ROM/RA3 ),
    .I1(\PCI-ROM/RB3 ),
    .I2(\PCI-ROM/RE3 ),
    .I3(\PCI-ROM/ROM3 ),
    .O(MD3)
  );
  X_OR4   \PCI-ROM/$1I8589  (
    .I0(\PCI-ROM/RA4 ),
    .I1(\PCI-ROM/RB4 ),
    .I2(\PCI-ROM/RE4 ),
    .I3(\PCI-ROM/ROM4 ),
    .O(MD4)
  );
  X_OR4   \PCI-ROM/$1I8588  (
    .I0(\PCI-ROM/RA5 ),
    .I1(\PCI-ROM/RB5 ),
    .I2(\PCI-ROM/RE5 ),
    .I3(\PCI-ROM/ROM5 ),
    .O(MD5)
  );
  X_OR4   \PCI-ROM/$1I8587  (
    .I0(\PCI-ROM/RA6 ),
    .I1(\PCI-ROM/RB6 ),
    .I2(\PCI-ROM/RE6 ),
    .I3(\PCI-ROM/ROM6 ),
    .O(MD6)
  );
  X_OR4   \PCI-ROM/$1I8586  (
    .I0(\PCI-ROM/RA7 ),
    .I1(\PCI-ROM/RB7 ),
    .I2(\PCI-ROM/RE7 ),
    .I3(\PCI-ROM/ROM7 ),
    .O(MD7)
  );
  X_OR4   \PCI-ROM/$1I8585  (
    .I0(\PCI-ROM/RA8 ),
    .I1(\PCI-ROM/RB8 ),
    .I2(\PCI-ROM/RE8 ),
    .I3(\PCI-ROM/ROM8 ),
    .O(MD8)
  );
  X_OR4   \PCI-ROM/$1I8584  (
    .I0(\PCI-ROM/RA9 ),
    .I1(\PCI-ROM/RB9 ),
    .I2(\PCI-ROM/RE9 ),
    .I3(\PCI-ROM/ROM9 ),
    .O(MD9)
  );
  X_OR4   \PCI-ROM/$1I8583  (
    .I0(\PCI-ROM/RA10 ),
    .I1(\PCI-ROM/RB10 ),
    .I2(\PCI-ROM/RE10 ),
    .I3(\PCI-ROM/ROM10 ),
    .O(MD10)
  );
  X_OR4   \PCI-ROM/$1I8582  (
    .I0(\PCI-ROM/RA11 ),
    .I1(\PCI-ROM/RB11 ),
    .I2(\PCI-ROM/RE11 ),
    .I3(\PCI-ROM/ROM11 ),
    .O(MD11)
  );
  X_OR4   \PCI-ROM/$1I8581  (
    .I0(\PCI-ROM/RA12 ),
    .I1(\PCI-ROM/RB12 ),
    .I2(\PCI-ROM/RE12 ),
    .I3(\PCI-ROM/ROM12 ),
    .O(MD12)
  );
  X_OR4   \PCI-ROM/$1I8580  (
    .I0(\PCI-ROM/RA13 ),
    .I1(\PCI-ROM/RB13 ),
    .I2(\PCI-ROM/RE13 ),
    .I3(\PCI-ROM/ROM13 ),
    .O(MD13)
  );
  X_OR4   \PCI-ROM/$1I8579  (
    .I0(\PCI-ROM/RA14 ),
    .I1(\PCI-ROM/RB14 ),
    .I2(\PCI-ROM/RE14 ),
    .I3(\PCI-ROM/ROM14 ),
    .O(MD14)
  );
  X_OR4   \PCI-ROM/$1I8578  (
    .I0(\PCI-ROM/RA15 ),
    .I1(\PCI-ROM/RB15 ),
    .I2(\PCI-ROM/RE15 ),
    .I3(\PCI-ROM/ROM15 ),
    .O(MD15)
  );
  X_OR4   \PCI-ROM/$1I8577  (
    .I0(\PCI-ROM/RA16 ),
    .I1(\PCI-ROM/RB16 ),
    .I2(\PCI-ROM/RE16 ),
    .I3(\PCI-ROM/ROM16 ),
    .O(MD16)
  );
  X_OR4   \PCI-ROM/$1I8576  (
    .I0(\PCI-ROM/RA17 ),
    .I1(\PCI-ROM/RB17 ),
    .I2(\PCI-ROM/RE17 ),
    .I3(\PCI-ROM/ROM17 ),
    .O(MD17)
  );
  X_OR4   \PCI-ROM/$1I8575  (
    .I0(\PCI-ROM/RA18 ),
    .I1(\PCI-ROM/RB18 ),
    .I2(\PCI-ROM/RE18 ),
    .I3(\PCI-ROM/ROM18 ),
    .O(MD18)
  );
  X_OR4   \PCI-ROM/$1I8574  (
    .I0(\PCI-ROM/RA19 ),
    .I1(\PCI-ROM/RB19 ),
    .I2(\PCI-ROM/RE19 ),
    .I3(\PCI-ROM/ROM19 ),
    .O(MD19)
  );
  X_OR4   \PCI-ROM/$1I8573  (
    .I0(\PCI-ROM/RA20 ),
    .I1(\PCI-ROM/RB20 ),
    .I2(\PCI-ROM/RE20 ),
    .I3(\PCI-ROM/ROM20 ),
    .O(MD20)
  );
  X_OR4   \PCI-ROM/$1I8572  (
    .I0(\PCI-ROM/RA21 ),
    .I1(\PCI-ROM/RB21 ),
    .I2(\PCI-ROM/RE21 ),
    .I3(\PCI-ROM/ROM21 ),
    .O(MD21)
  );
  X_OR4   \PCI-ROM/$1I8571  (
    .I0(\PCI-ROM/RA22 ),
    .I1(\PCI-ROM/RB22 ),
    .I2(\PCI-ROM/RE22 ),
    .I3(\PCI-ROM/ROM22 ),
    .O(MD22)
  );
  X_OR4   \PCI-ROM/$1I8570  (
    .I0(\PCI-ROM/RA23 ),
    .I1(\PCI-ROM/RB23 ),
    .I2(\PCI-ROM/RE23 ),
    .I3(\PCI-ROM/ROM23 ),
    .O(MD23)
  );
  X_OR4   \PCI-ROM/$1I8569  (
    .I0(\PCI-ROM/RA24 ),
    .I1(\PCI-ROM/RB24 ),
    .I2(\PCI-ROM/RE24 ),
    .I3(\PCI-ROM/ROM24 ),
    .O(MD24)
  );
  X_OR4   \PCI-ROM/$1I8568  (
    .I0(\PCI-ROM/RA25 ),
    .I1(\PCI-ROM/RB25 ),
    .I2(\PCI-ROM/RE25 ),
    .I3(\PCI-ROM/ROM25 ),
    .O(MD25)
  );
  X_OR4   \PCI-ROM/$1I8567  (
    .I0(\PCI-ROM/RA26 ),
    .I1(\PCI-ROM/RB26 ),
    .I2(\PCI-ROM/RE26 ),
    .I3(\PCI-ROM/ROM26 ),
    .O(MD26)
  );
  X_OR4   \PCI-ROM/$1I8566  (
    .I0(\PCI-ROM/RA27 ),
    .I1(\PCI-ROM/RB27 ),
    .I2(\PCI-ROM/RE27 ),
    .I3(\PCI-ROM/ROM27 ),
    .O(MD27)
  );
  X_OR4   \PCI-ROM/$1I8565  (
    .I0(\PCI-ROM/RA28 ),
    .I1(\PCI-ROM/RB28 ),
    .I2(\PCI-ROM/RE28 ),
    .I3(\PCI-ROM/ROM28 ),
    .O(MD28)
  );
  X_OR4   \PCI-ROM/$1I8564  (
    .I0(\PCI-ROM/RA29 ),
    .I1(\PCI-ROM/RB29 ),
    .I2(\PCI-ROM/RE29 ),
    .I3(\PCI-ROM/ROM29 ),
    .O(MD29)
  );
  X_OR4   \PCI-ROM/$1I8563  (
    .I0(\PCI-ROM/RA30 ),
    .I1(\PCI-ROM/RB30 ),
    .I2(\PCI-ROM/RE30 ),
    .I3(\PCI-ROM/ROM30 ),
    .O(MD30)
  );
  X_OR4   \PCI-ROM/$1I8562  (
    .I0(\PCI-ROM/RA31 ),
    .I1(\PCI-ROM/RB31 ),
    .I2(\PCI-ROM/RE31 ),
    .I3(\PCI-ROM/ROM31 ),
    .O(MD31)
  );
  X_OR3   \PCI-ROM/$1I8561  (
    .I0(\PCI-ROM/RC0 ),
    .I1(\PCI-ROM/RF0 ),
    .I2(\PCI-ROM/RD0 ),
    .O(\PCI-ROM/ROM0 )
  );
  X_OR3   \PCI-ROM/$1I8560  (
    .I0(\PCI-ROM/RC1 ),
    .I1(\PCI-ROM/RF1 ),
    .I2(\PCI-ROM/RD1 ),
    .O(\PCI-ROM/ROM1 )
  );
  X_OR3   \PCI-ROM/$1I8559  (
    .I0(\PCI-ROM/RC2 ),
    .I1(\PCI-ROM/RF2 ),
    .I2(\PCI-ROM/RD2 ),
    .O(\PCI-ROM/ROM2 )
  );
  X_OR3   \PCI-ROM/$1I8558  (
    .I0(\PCI-ROM/RC3 ),
    .I1(\PCI-ROM/RF3 ),
    .I2(\PCI-ROM/RD3 ),
    .O(\PCI-ROM/ROM3 )
  );
  X_OR3   \PCI-ROM/$1I8557  (
    .I0(\PCI-ROM/RC4 ),
    .I1(\PCI-ROM/RF4 ),
    .I2(\PCI-ROM/RD4 ),
    .O(\PCI-ROM/ROM4 )
  );
  X_OR3   \PCI-ROM/$1I8556  (
    .I0(\PCI-ROM/RC5 ),
    .I1(\PCI-ROM/RF5 ),
    .I2(\PCI-ROM/RD5 ),
    .O(\PCI-ROM/ROM5 )
  );
  X_OR3   \PCI-ROM/$1I8555  (
    .I0(\PCI-ROM/RC6 ),
    .I1(\PCI-ROM/RF6 ),
    .I2(\PCI-ROM/RD6 ),
    .O(\PCI-ROM/ROM6 )
  );
  X_OR3   \PCI-ROM/$1I8554  (
    .I0(\PCI-ROM/RC7 ),
    .I1(\PCI-ROM/RF7 ),
    .I2(\PCI-ROM/RD7 ),
    .O(\PCI-ROM/ROM7 )
  );
  X_OR3   \PCI-ROM/$1I8553  (
    .I0(\PCI-ROM/RC8 ),
    .I1(\PCI-ROM/RF8 ),
    .I2(\PCI-ROM/RD8 ),
    .O(\PCI-ROM/ROM8 )
  );
  X_OR3   \PCI-ROM/$1I8552  (
    .I0(\PCI-ROM/RC9 ),
    .I1(\PCI-ROM/RF9 ),
    .I2(\PCI-ROM/RD9 ),
    .O(\PCI-ROM/ROM9 )
  );
  X_OR3   \PCI-ROM/$1I8551  (
    .I0(\PCI-ROM/RC10 ),
    .I1(\PCI-ROM/RF10 ),
    .I2(\PCI-ROM/RD10 ),
    .O(\PCI-ROM/ROM10 )
  );
  X_OR3   \PCI-ROM/$1I8550  (
    .I0(\PCI-ROM/RC11 ),
    .I1(\PCI-ROM/RF11 ),
    .I2(\PCI-ROM/RD11 ),
    .O(\PCI-ROM/ROM11 )
  );
  X_OR3   \PCI-ROM/$1I8549  (
    .I0(\PCI-ROM/RC12 ),
    .I1(\PCI-ROM/RF12 ),
    .I2(\PCI-ROM/RD12 ),
    .O(\PCI-ROM/ROM12 )
  );
  X_OR3   \PCI-ROM/$1I8548  (
    .I0(\PCI-ROM/RC13 ),
    .I1(\PCI-ROM/RF13 ),
    .I2(\PCI-ROM/RD13 ),
    .O(\PCI-ROM/ROM13 )
  );
  X_OR3   \PCI-ROM/$1I8547  (
    .I0(\PCI-ROM/RC14 ),
    .I1(\PCI-ROM/RF14 ),
    .I2(\PCI-ROM/RD14 ),
    .O(\PCI-ROM/ROM14 )
  );
  X_OR3   \PCI-ROM/$1I8546  (
    .I0(\PCI-ROM/RC15 ),
    .I1(\PCI-ROM/RF15 ),
    .I2(\PCI-ROM/RD15 ),
    .O(\PCI-ROM/ROM15 )
  );
  X_OR3   \PCI-ROM/$1I8545  (
    .I0(\PCI-ROM/RC16 ),
    .I1(\PCI-ROM/RF16 ),
    .I2(\PCI-ROM/RD16 ),
    .O(\PCI-ROM/ROM16 )
  );
  X_OR3   \PCI-ROM/$1I8544  (
    .I0(\PCI-ROM/RC17 ),
    .I1(\PCI-ROM/RF17 ),
    .I2(\PCI-ROM/RD17 ),
    .O(\PCI-ROM/ROM17 )
  );
  X_OR3   \PCI-ROM/$1I8543  (
    .I0(\PCI-ROM/RC18 ),
    .I1(\PCI-ROM/RF18 ),
    .I2(\PCI-ROM/RD18 ),
    .O(\PCI-ROM/ROM18 )
  );
  X_OR3   \PCI-ROM/$1I8542  (
    .I0(\PCI-ROM/RC19 ),
    .I1(\PCI-ROM/RF19 ),
    .I2(\PCI-ROM/RD19 ),
    .O(\PCI-ROM/ROM19 )
  );
  X_OR3   \PCI-ROM/$1I8541  (
    .I0(\PCI-ROM/RC20 ),
    .I1(\PCI-ROM/RF20 ),
    .I2(\PCI-ROM/RD20 ),
    .O(\PCI-ROM/ROM20 )
  );
  X_OR3   \PCI-ROM/$1I8540  (
    .I0(\PCI-ROM/RC21 ),
    .I1(\PCI-ROM/RF21 ),
    .I2(\PCI-ROM/RD21 ),
    .O(\PCI-ROM/ROM21 )
  );
  X_OR3   \PCI-ROM/$1I8539  (
    .I0(\PCI-ROM/RC22 ),
    .I1(\PCI-ROM/RF22 ),
    .I2(\PCI-ROM/RD22 ),
    .O(\PCI-ROM/ROM22 )
  );
  X_OR3   \PCI-ROM/$1I8538  (
    .I0(\PCI-ROM/RC23 ),
    .I1(\PCI-ROM/RF23 ),
    .I2(\PCI-ROM/RD23 ),
    .O(\PCI-ROM/ROM23 )
  );
  X_OR3   \PCI-ROM/$1I8537  (
    .I0(\PCI-ROM/RC24 ),
    .I1(\PCI-ROM/RF24 ),
    .I2(\PCI-ROM/RD24 ),
    .O(\PCI-ROM/ROM24 )
  );
  X_OR3   \PCI-ROM/$1I8536  (
    .I0(\PCI-ROM/RC25 ),
    .I1(\PCI-ROM/RF25 ),
    .I2(\PCI-ROM/RD25 ),
    .O(\PCI-ROM/ROM25 )
  );
  X_OR3   \PCI-ROM/$1I8535  (
    .I0(\PCI-ROM/RC26 ),
    .I1(\PCI-ROM/RF26 ),
    .I2(\PCI-ROM/RD26 ),
    .O(\PCI-ROM/ROM26 )
  );
  X_OR3   \PCI-ROM/$1I8534  (
    .I0(\PCI-ROM/RC27 ),
    .I1(\PCI-ROM/RF27 ),
    .I2(\PCI-ROM/RD27 ),
    .O(\PCI-ROM/ROM27 )
  );
  X_OR3   \PCI-ROM/$1I8533  (
    .I0(\PCI-ROM/RC28 ),
    .I1(\PCI-ROM/RF28 ),
    .I2(\PCI-ROM/RD28 ),
    .O(\PCI-ROM/ROM28 )
  );
  X_OR3   \PCI-ROM/$1I8532  (
    .I0(\PCI-ROM/RC29 ),
    .I1(\PCI-ROM/RF29 ),
    .I2(\PCI-ROM/RD29 ),
    .O(\PCI-ROM/ROM29 )
  );
  X_OR3   \PCI-ROM/$1I8531  (
    .I0(\PCI-ROM/RC30 ),
    .I1(\PCI-ROM/RF30 ),
    .I2(\PCI-ROM/RD30 ),
    .O(\PCI-ROM/ROM30 )
  );
  X_OR3   \PCI-ROM/$1I8530  (
    .I0(\PCI-ROM/RC31 ),
    .I1(\PCI-ROM/RF31 ),
    .I2(\PCI-ROM/RD31 ),
    .O(\PCI-ROM/ROM31 )
  );
  X_BUF   \PCI-ROM/$1I8478  (
    .I(\PCI-ROM/$1N8453 ),
    .O(\PCI-ROM/CLR8 )
  );
  X_BUF   \PCI-ROM/$1I8477  (
    .I(\PCI-ROM/$1N8453 ),
    .O(\PCI-ROM/CLR9 )
  );
  X_BUF   \PCI-ROM/$1I8476  (
    .I(\PCI-ROM/$1N8453 ),
    .O(\PCI-ROM/CLR10 )
  );
  X_BUF   \PCI-ROM/$1I8475  (
    .I(\PCI-ROM/$1N8453 ),
    .O(\PCI-ROM/CLR11 )
  );
  X_BUF   \PCI-ROM/$1I8474  (
    .I(\PCI-ROM/$1N8453 ),
    .O(\PCI-ROM/CLR12 )
  );
  X_BUF   \PCI-ROM/$1I8473  (
    .I(\PCI-ROM/$1N8453 ),
    .O(\PCI-ROM/CLR13 )
  );
  X_BUF   \PCI-ROM/$1I8472  (
    .I(\PCI-ROM/$1N8453 ),
    .O(\PCI-ROM/CLR14 )
  );
  X_BUF   \PCI-ROM/$1I8471  (
    .I(\PCI-ROM/$1N8453 ),
    .O(\PCI-ROM/CLR15 )
  );
  X_BUF   \PCI-ROM/$1I8470  (
    .I(\PCI-ROM/$1N8453 ),
    .O(\PCI-ROM/CLR16 )
  );
  X_BUF   \PCI-ROM/$1I8469  (
    .I(\PCI-ROM/$1N8453 ),
    .O(\PCI-ROM/CLR17 )
  );
  X_BUF   \PCI-ROM/$1I8468  (
    .I(\PCI-ROM/$1N8453 ),
    .O(\PCI-ROM/CLR18 )
  );
  X_BUF   \PCI-ROM/$1I8467  (
    .I(\PCI-ROM/$1N8453 ),
    .O(\PCI-ROM/CLR19 )
  );
  X_BUF   \PCI-ROM/$1I8466  (
    .I(\PCI-ROM/$1N8453 ),
    .O(\PCI-ROM/CLR20 )
  );
  X_BUF   \PCI-ROM/$1I8465  (
    .I(\PCI-ROM/$1N8453 ),
    .O(\PCI-ROM/CLR21 )
  );
  X_BUF   \PCI-ROM/$1I8464  (
    .I(\PCI-ROM/$1N8453 ),
    .O(\PCI-ROM/CLR22 )
  );
  X_BUF   \PCI-ROM/$1I8463  (
    .I(\PCI-ROM/$1N8453 ),
    .O(\PCI-ROM/CLR23 )
  );
  X_BUF   \PCI-ROM/$1I8462  (
    .I(\PCI-ROM/$1N8453 ),
    .O(\PCI-ROM/CLR24 )
  );
  X_BUF   \PCI-ROM/$1I8461  (
    .I(\PCI-ROM/$1N8453 ),
    .O(\PCI-ROM/CLR25 )
  );
  X_BUF   \PCI-ROM/$1I8460  (
    .I(\PCI-ROM/$1N8453 ),
    .O(\PCI-ROM/CLR26 )
  );
  X_BUF   \PCI-ROM/$1I8459  (
    .I(\PCI-ROM/$1N8453 ),
    .O(\PCI-ROM/CLR27 )
  );
  X_BUF   \PCI-ROM/$1I8458  (
    .I(\PCI-ROM/$1N8453 ),
    .O(\PCI-ROM/CLR28 )
  );
  X_BUF   \PCI-ROM/$1I8457  (
    .I(\PCI-ROM/$1N8453 ),
    .O(\PCI-ROM/CLR29 )
  );
  X_BUF   \PCI-ROM/$1I8456  (
    .I(\PCI-ROM/$1N8453 ),
    .O(\PCI-ROM/CLR30 )
  );
  X_BUF   \PCI-ROM/$1I8455  (
    .I(\PCI-ROM/$1N8453 ),
    .O(\PCI-ROM/CLR31 )
  );
  X_BUF   \PCI-ROM/$1I8434  (
    .I(CFG232),
    .O(\PCI-ROM/CLR0 )
  );
  X_BUF   \PCI-ROM/$1I8433  (
    .I(CFG233),
    .O(\PCI-ROM/CLR1 )
  );
  X_BUF   \PCI-ROM/$1I8432  (
    .I(CFG234),
    .O(\PCI-ROM/CLR2 )
  );
  X_BUF   \PCI-ROM/$1I8431  (
    .I(CFG235),
    .O(\PCI-ROM/CLR3 )
  );
  X_BUF   \PCI-ROM/$1I8430  (
    .I(CFG236),
    .O(\PCI-ROM/CLR4 )
  );
  X_BUF   \PCI-ROM/$1I8429  (
    .I(CFG237),
    .O(\PCI-ROM/CLR5 )
  );
  X_BUF   \PCI-ROM/$1I8428  (
    .I(CFG238),
    .O(\PCI-ROM/CLR6 )
  );
  X_BUF   \PCI-ROM/$1I8427  (
    .I(CFG239),
    .O(\PCI-ROM/CLR7 )
  );
  X_AND2   \PCI-ROM/$1I8365  (
    .I0(\PCI-ROM/SELD ),
    .I1(\PCI-ROM/CLR0 ),
    .O(\PCI-ROM/RF0 )
  );
  X_AND2   \PCI-ROM/$1I8364  (
    .I0(\PCI-ROM/SELD ),
    .I1(\PCI-ROM/CLR1 ),
    .O(\PCI-ROM/RF1 )
  );
  X_AND2   \PCI-ROM/$1I8363  (
    .I0(\PCI-ROM/SELD ),
    .I1(\PCI-ROM/CLR2 ),
    .O(\PCI-ROM/RF2 )
  );
  X_AND2   \PCI-ROM/$1I8362  (
    .I0(\PCI-ROM/SELD ),
    .I1(\PCI-ROM/CLR3 ),
    .O(\PCI-ROM/RF3 )
  );
  X_AND2   \PCI-ROM/$1I8361  (
    .I0(\PCI-ROM/SELD ),
    .I1(\PCI-ROM/CLR4 ),
    .O(\PCI-ROM/RF4 )
  );
  X_AND2   \PCI-ROM/$1I8360  (
    .I0(\PCI-ROM/SELD ),
    .I1(\PCI-ROM/CLR5 ),
    .O(\PCI-ROM/RF5 )
  );
  X_AND2   \PCI-ROM/$1I8359  (
    .I0(\PCI-ROM/SELD ),
    .I1(\PCI-ROM/CLR6 ),
    .O(\PCI-ROM/RF6 )
  );
  X_AND2   \PCI-ROM/$1I8358  (
    .I0(\PCI-ROM/SELD ),
    .I1(\PCI-ROM/CLR7 ),
    .O(\PCI-ROM/RF7 )
  );
  X_AND2   \PCI-ROM/$1I8357  (
    .I0(\PCI-ROM/SELD ),
    .I1(\PCI-ROM/CLR8 ),
    .O(\PCI-ROM/RF8 )
  );
  X_AND2   \PCI-ROM/$1I8356  (
    .I0(\PCI-ROM/SELD ),
    .I1(\PCI-ROM/CLR9 ),
    .O(\PCI-ROM/RF9 )
  );
  X_AND2   \PCI-ROM/$1I8355  (
    .I0(\PCI-ROM/SELD ),
    .I1(\PCI-ROM/CLR10 ),
    .O(\PCI-ROM/RF10 )
  );
  X_AND2   \PCI-ROM/$1I8354  (
    .I0(\PCI-ROM/SELD ),
    .I1(\PCI-ROM/CLR11 ),
    .O(\PCI-ROM/RF11 )
  );
  X_AND2   \PCI-ROM/$1I8353  (
    .I0(\PCI-ROM/SELD ),
    .I1(\PCI-ROM/CLR12 ),
    .O(\PCI-ROM/RF12 )
  );
  X_AND2   \PCI-ROM/$1I8352  (
    .I0(\PCI-ROM/SELD ),
    .I1(\PCI-ROM/CLR13 ),
    .O(\PCI-ROM/RF13 )
  );
  X_AND2   \PCI-ROM/$1I8351  (
    .I0(\PCI-ROM/SELD ),
    .I1(\PCI-ROM/CLR14 ),
    .O(\PCI-ROM/RF14 )
  );
  X_AND2   \PCI-ROM/$1I8350  (
    .I0(\PCI-ROM/SELD ),
    .I1(\PCI-ROM/CLR15 ),
    .O(\PCI-ROM/RF15 )
  );
  X_AND2   \PCI-ROM/$1I8349  (
    .I0(\PCI-ROM/SELD ),
    .I1(\PCI-ROM/CLR16 ),
    .O(\PCI-ROM/RF16 )
  );
  X_AND2   \PCI-ROM/$1I8348  (
    .I0(\PCI-ROM/SELD ),
    .I1(\PCI-ROM/CLR17 ),
    .O(\PCI-ROM/RF17 )
  );
  X_AND2   \PCI-ROM/$1I8347  (
    .I0(\PCI-ROM/SELD ),
    .I1(\PCI-ROM/CLR18 ),
    .O(\PCI-ROM/RF18 )
  );
  X_AND2   \PCI-ROM/$1I8346  (
    .I0(\PCI-ROM/SELD ),
    .I1(\PCI-ROM/CLR19 ),
    .O(\PCI-ROM/RF19 )
  );
  X_AND2   \PCI-ROM/$1I8345  (
    .I0(\PCI-ROM/SELD ),
    .I1(\PCI-ROM/CLR20 ),
    .O(\PCI-ROM/RF20 )
  );
  X_AND2   \PCI-ROM/$1I8344  (
    .I0(\PCI-ROM/SELD ),
    .I1(\PCI-ROM/CLR21 ),
    .O(\PCI-ROM/RF21 )
  );
  X_AND2   \PCI-ROM/$1I8343  (
    .I0(\PCI-ROM/SELD ),
    .I1(\PCI-ROM/CLR22 ),
    .O(\PCI-ROM/RF22 )
  );
  X_AND2   \PCI-ROM/$1I8342  (
    .I0(\PCI-ROM/SELD ),
    .I1(\PCI-ROM/CLR23 ),
    .O(\PCI-ROM/RF23 )
  );
  X_AND2   \PCI-ROM/$1I8341  (
    .I0(\PCI-ROM/SELD ),
    .I1(\PCI-ROM/CLR24 ),
    .O(\PCI-ROM/RF24 )
  );
  X_AND2   \PCI-ROM/$1I8340  (
    .I0(\PCI-ROM/SELD ),
    .I1(\PCI-ROM/CLR25 ),
    .O(\PCI-ROM/RF25 )
  );
  X_AND2   \PCI-ROM/$1I8339  (
    .I0(\PCI-ROM/SELD ),
    .I1(\PCI-ROM/CLR26 ),
    .O(\PCI-ROM/RF26 )
  );
  X_AND2   \PCI-ROM/$1I8338  (
    .I0(\PCI-ROM/SELD ),
    .I1(\PCI-ROM/CLR27 ),
    .O(\PCI-ROM/RF27 )
  );
  X_AND2   \PCI-ROM/$1I8337  (
    .I0(\PCI-ROM/SELD ),
    .I1(\PCI-ROM/CLR28 ),
    .O(\PCI-ROM/RF28 )
  );
  X_AND2   \PCI-ROM/$1I8336  (
    .I0(\PCI-ROM/SELD ),
    .I1(\PCI-ROM/CLR29 ),
    .O(\PCI-ROM/RF29 )
  );
  X_AND2   \PCI-ROM/$1I8335  (
    .I0(\PCI-ROM/SELD ),
    .I1(\PCI-ROM/CLR30 ),
    .O(\PCI-ROM/RF30 )
  );
  X_AND2   \PCI-ROM/$1I8334  (
    .I0(\PCI-ROM/SELD ),
    .I1(\PCI-ROM/CLR31 ),
    .O(\PCI-ROM/RF31 )
  );
  X_AND4   \PCI-ROM/$1I8330  (
    .I0(\NlwInverterSignal_PCI-ROM/$1I8330/I0 ),
    .I1(\NlwInverterSignal_PCI-ROM/$1I8330/I1 ),
    .I2(CFG116),
    .I3(\PCI-ROM/$1N8328 ),
    .O(\PCI-ROM/SELD )
  );
  X_AND2   \PCI-ROM/$1I8321  (
    .I0(\PCI-ROM/SELBY ),
    .I1(CFG184),
    .O(\PCI-ROM/RE0 )
  );
  X_AND2   \PCI-ROM/$1I8320  (
    .I0(\PCI-ROM/SELBY ),
    .I1(CFG185),
    .O(\PCI-ROM/RE1 )
  );
  X_AND2   \PCI-ROM/$1I8319  (
    .I0(\PCI-ROM/SELBY ),
    .I1(CFG186),
    .O(\PCI-ROM/RE2 )
  );
  X_AND2   \PCI-ROM/$1I8318  (
    .I0(\PCI-ROM/SELBY ),
    .I1(CFG187),
    .O(\PCI-ROM/RE3 )
  );
  X_AND2   \PCI-ROM/$1I8317  (
    .I0(\PCI-ROM/SELBY ),
    .I1(CFG188),
    .O(\PCI-ROM/RE4 )
  );
  X_AND2   \PCI-ROM/$1I8316  (
    .I0(\PCI-ROM/SELBY ),
    .I1(CFG189),
    .O(\PCI-ROM/RE5 )
  );
  X_AND2   \PCI-ROM/$1I8315  (
    .I0(\PCI-ROM/SELBY ),
    .I1(CFG190),
    .O(\PCI-ROM/RE6 )
  );
  X_AND2   \PCI-ROM/$1I8314  (
    .I0(\PCI-ROM/SELBY ),
    .I1(CFG191),
    .O(\PCI-ROM/RE7 )
  );
  X_AND2   \PCI-ROM/$1I8313  (
    .I0(\PCI-ROM/SELBY ),
    .I1(CFG192),
    .O(\PCI-ROM/RE8 )
  );
  X_AND2   \PCI-ROM/$1I8312  (
    .I0(\PCI-ROM/SELBY ),
    .I1(CFG193),
    .O(\PCI-ROM/RE9 )
  );
  X_AND2   \PCI-ROM/$1I8311  (
    .I0(\PCI-ROM/SELBY ),
    .I1(CFG194),
    .O(\PCI-ROM/RE10 )
  );
  X_AND2   \PCI-ROM/$1I8310  (
    .I0(\PCI-ROM/SELBY ),
    .I1(CFG195),
    .O(\PCI-ROM/RE11 )
  );
  X_AND2   \PCI-ROM/$1I8309  (
    .I0(\PCI-ROM/SELBY ),
    .I1(CFG196),
    .O(\PCI-ROM/RE12 )
  );
  X_AND2   \PCI-ROM/$1I8308  (
    .I0(\PCI-ROM/SELBY ),
    .I1(CFG197),
    .O(\PCI-ROM/RE13 )
  );
  X_AND2   \PCI-ROM/$1I8307  (
    .I0(\PCI-ROM/SELBY ),
    .I1(CFG198),
    .O(\PCI-ROM/RE14 )
  );
  X_AND2   \PCI-ROM/$1I8306  (
    .I0(\PCI-ROM/SELBY ),
    .I1(CFG199),
    .O(\PCI-ROM/RE15 )
  );
  X_AND2   \PCI-ROM/$1I8305  (
    .I0(\PCI-ROM/SELBY ),
    .I1(CFG200),
    .O(\PCI-ROM/RE16 )
  );
  X_AND2   \PCI-ROM/$1I8304  (
    .I0(\PCI-ROM/SELBY ),
    .I1(CFG201),
    .O(\PCI-ROM/RE17 )
  );
  X_AND2   \PCI-ROM/$1I8303  (
    .I0(\PCI-ROM/SELBY ),
    .I1(CFG202),
    .O(\PCI-ROM/RE18 )
  );
  X_AND2   \PCI-ROM/$1I8302  (
    .I0(\PCI-ROM/SELBY ),
    .I1(CFG203),
    .O(\PCI-ROM/RE19 )
  );
  X_AND2   \PCI-ROM/$1I8301  (
    .I0(\PCI-ROM/SELBY ),
    .I1(CFG204),
    .O(\PCI-ROM/RE20 )
  );
  X_AND2   \PCI-ROM/$1I8300  (
    .I0(\PCI-ROM/SELBY ),
    .I1(CFG205),
    .O(\PCI-ROM/RE21 )
  );
  X_AND2   \PCI-ROM/$1I8299  (
    .I0(\PCI-ROM/SELBY ),
    .I1(CFG206),
    .O(\PCI-ROM/RE22 )
  );
  X_AND2   \PCI-ROM/$1I8298  (
    .I0(\PCI-ROM/SELBY ),
    .I1(CFG207),
    .O(\PCI-ROM/RE23 )
  );
  X_AND2   \PCI-ROM/$1I8297  (
    .I0(\PCI-ROM/SELBY ),
    .I1(CFG208),
    .O(\PCI-ROM/RE24 )
  );
  X_AND2   \PCI-ROM/$1I8296  (
    .I0(\PCI-ROM/SELBY ),
    .I1(CFG209),
    .O(\PCI-ROM/RE25 )
  );
  X_AND2   \PCI-ROM/$1I8295  (
    .I0(\PCI-ROM/SELBY ),
    .I1(CFG210),
    .O(\PCI-ROM/RE26 )
  );
  X_AND2   \PCI-ROM/$1I8294  (
    .I0(\PCI-ROM/SELBY ),
    .I1(CFG211),
    .O(\PCI-ROM/RE27 )
  );
  X_AND2   \PCI-ROM/$1I8293  (
    .I0(\PCI-ROM/SELBY ),
    .I1(CFG212),
    .O(\PCI-ROM/RE28 )
  );
  X_AND2   \PCI-ROM/$1I8292  (
    .I0(\PCI-ROM/SELBY ),
    .I1(CFG213),
    .O(\PCI-ROM/RE29 )
  );
  X_AND2   \PCI-ROM/$1I8291  (
    .I0(\PCI-ROM/SELBY ),
    .I1(CFG214),
    .O(\PCI-ROM/RE30 )
  );
  X_AND2   \PCI-ROM/$1I8290  (
    .I0(\PCI-ROM/SELBY ),
    .I1(CFG215),
    .O(\PCI-ROM/RE31 )
  );
  X_AND4   \PCI-ROM/$1I8282  (
    .I0(\NlwInverterSignal_PCI-ROM/$1I8282/I0 ),
    .I1(\NlwInverterSignal_PCI-ROM/$1I8282/I1 ),
    .I2(\NlwInverterSignal_PCI-ROM/$1I8282/I2 ),
    .I3(\PCI-ROM/$1N8283 ),
    .O(\PCI-ROM/SELBY )
  );
  X_AND2   \PCI-ROM/$1I8275  (
    .I0(\PCI-ROM/SELBX ),
    .I1(SUB_DATA0),
    .O(\PCI-ROM/RD0 )
  );
  X_AND2   \PCI-ROM/$1I8274  (
    .I0(\PCI-ROM/SELBX ),
    .I1(SUB_DATA1),
    .O(\PCI-ROM/RD1 )
  );
  X_AND2   \PCI-ROM/$1I8273  (
    .I0(\PCI-ROM/SELBX ),
    .I1(SUB_DATA2),
    .O(\PCI-ROM/RD2 )
  );
  X_AND2   \PCI-ROM/$1I8272  (
    .I0(\PCI-ROM/SELBX ),
    .I1(SUB_DATA3),
    .O(\PCI-ROM/RD3 )
  );
  X_AND2   \PCI-ROM/$1I8271  (
    .I0(\PCI-ROM/SELBX ),
    .I1(SUB_DATA4),
    .O(\PCI-ROM/RD4 )
  );
  X_AND2   \PCI-ROM/$1I8270  (
    .I0(\PCI-ROM/SELBX ),
    .I1(SUB_DATA5),
    .O(\PCI-ROM/RD5 )
  );
  X_AND2   \PCI-ROM/$1I8269  (
    .I0(\PCI-ROM/SELBX ),
    .I1(SUB_DATA6),
    .O(\PCI-ROM/RD6 )
  );
  X_AND2   \PCI-ROM/$1I8268  (
    .I0(\PCI-ROM/SELBX ),
    .I1(SUB_DATA7),
    .O(\PCI-ROM/RD7 )
  );
  X_AND2   \PCI-ROM/$1I8267  (
    .I0(\PCI-ROM/SELBX ),
    .I1(SUB_DATA8),
    .O(\PCI-ROM/RD8 )
  );
  X_AND2   \PCI-ROM/$1I8266  (
    .I0(\PCI-ROM/SELBX ),
    .I1(SUB_DATA9),
    .O(\PCI-ROM/RD9 )
  );
  X_AND2   \PCI-ROM/$1I8265  (
    .I0(\PCI-ROM/SELBX ),
    .I1(SUB_DATA10),
    .O(\PCI-ROM/RD10 )
  );
  X_AND2   \PCI-ROM/$1I8264  (
    .I0(\PCI-ROM/SELBX ),
    .I1(SUB_DATA11),
    .O(\PCI-ROM/RD11 )
  );
  X_AND2   \PCI-ROM/$1I8263  (
    .I0(\PCI-ROM/SELBX ),
    .I1(SUB_DATA12),
    .O(\PCI-ROM/RD12 )
  );
  X_AND2   \PCI-ROM/$1I8262  (
    .I0(\PCI-ROM/SELBX ),
    .I1(SUB_DATA13),
    .O(\PCI-ROM/RD13 )
  );
  X_AND2   \PCI-ROM/$1I8261  (
    .I0(\PCI-ROM/SELBX ),
    .I1(SUB_DATA14),
    .O(\PCI-ROM/RD14 )
  );
  X_AND2   \PCI-ROM/$1I8260  (
    .I0(\PCI-ROM/SELBX ),
    .I1(SUB_DATA15),
    .O(\PCI-ROM/RD15 )
  );
  X_AND2   \PCI-ROM/$1I8259  (
    .I0(\PCI-ROM/SELBX ),
    .I1(SUB_DATA16),
    .O(\PCI-ROM/RD16 )
  );
  X_AND2   \PCI-ROM/$1I8258  (
    .I0(\PCI-ROM/SELBX ),
    .I1(SUB_DATA17),
    .O(\PCI-ROM/RD17 )
  );
  X_AND2   \PCI-ROM/$1I8257  (
    .I0(\PCI-ROM/SELBX ),
    .I1(SUB_DATA18),
    .O(\PCI-ROM/RD18 )
  );
  X_AND2   \PCI-ROM/$1I8256  (
    .I0(\PCI-ROM/SELBX ),
    .I1(SUB_DATA19),
    .O(\PCI-ROM/RD19 )
  );
  X_AND2   \PCI-ROM/$1I8255  (
    .I0(\PCI-ROM/SELBX ),
    .I1(SUB_DATA20),
    .O(\PCI-ROM/RD20 )
  );
  X_AND2   \PCI-ROM/$1I8254  (
    .I0(\PCI-ROM/SELBX ),
    .I1(SUB_DATA21),
    .O(\PCI-ROM/RD21 )
  );
  X_AND2   \PCI-ROM/$1I8253  (
    .I0(\PCI-ROM/SELBX ),
    .I1(SUB_DATA22),
    .O(\PCI-ROM/RD22 )
  );
  X_AND2   \PCI-ROM/$1I8252  (
    .I0(\PCI-ROM/SELBX ),
    .I1(SUB_DATA23),
    .O(\PCI-ROM/RD23 )
  );
  X_AND2   \PCI-ROM/$1I8251  (
    .I0(\PCI-ROM/SELBX ),
    .I1(SUB_DATA24),
    .O(\PCI-ROM/RD24 )
  );
  X_AND2   \PCI-ROM/$1I8250  (
    .I0(\PCI-ROM/SELBX ),
    .I1(SUB_DATA25),
    .O(\PCI-ROM/RD25 )
  );
  X_AND2   \PCI-ROM/$1I8249  (
    .I0(\PCI-ROM/SELBX ),
    .I1(SUB_DATA26),
    .O(\PCI-ROM/RD26 )
  );
  X_AND2   \PCI-ROM/$1I8248  (
    .I0(\PCI-ROM/SELBX ),
    .I1(SUB_DATA27),
    .O(\PCI-ROM/RD27 )
  );
  X_AND2   \PCI-ROM/$1I8247  (
    .I0(\PCI-ROM/SELBX ),
    .I1(SUB_DATA28),
    .O(\PCI-ROM/RD28 )
  );
  X_AND2   \PCI-ROM/$1I8246  (
    .I0(\PCI-ROM/SELBX ),
    .I1(SUB_DATA29),
    .O(\PCI-ROM/RD29 )
  );
  X_AND2   \PCI-ROM/$1I8245  (
    .I0(\PCI-ROM/SELBX ),
    .I1(SUB_DATA30),
    .O(\PCI-ROM/RD30 )
  );
  X_AND2   \PCI-ROM/$1I8244  (
    .I0(\PCI-ROM/SELBX ),
    .I1(SUB_DATA31),
    .O(\PCI-ROM/RD31 )
  );
  X_AND4   \PCI-ROM/$1I8237  (
    .I0(\NlwInverterSignal_PCI-ROM/$1I8237/I0 ),
    .I1(\NlwInverterSignal_PCI-ROM/$1I8237/I1 ),
    .I2(CFG114),
    .I3(\PCI-ROM/$1N8238 ),
    .O(\PCI-ROM/SELBX )
  );
  X_AND4   \PCI-ROM/$1I8227  (
    .I0(\NlwInverterSignal_PCI-ROM/$1I8227/I0 ),
    .I1(\NlwInverterSignal_PCI-ROM/$1I8227/I1 ),
    .I2(\NlwInverterSignal_PCI-ROM/$1I8227/I2 ),
    .I3(\PCI-ROM/$1N8188 ),
    .O(\PCI-ROM/SELA )
  );
  X_AND2   \PCI-ROM/$1I8224  (
    .I0(\PCI-ROM/SELA ),
    .I1(SUB_DATA0),
    .O(\PCI-ROM/RC0 )
  );
  X_AND2   \PCI-ROM/$1I8223  (
    .I0(\PCI-ROM/SELA ),
    .I1(SUB_DATA1),
    .O(\PCI-ROM/RC1 )
  );
  X_AND2   \PCI-ROM/$1I8222  (
    .I0(\PCI-ROM/SELA ),
    .I1(SUB_DATA2),
    .O(\PCI-ROM/RC2 )
  );
  X_AND2   \PCI-ROM/$1I8221  (
    .I0(\PCI-ROM/SELA ),
    .I1(SUB_DATA3),
    .O(\PCI-ROM/RC3 )
  );
  X_AND2   \PCI-ROM/$1I8220  (
    .I0(\PCI-ROM/SELA ),
    .I1(SUB_DATA4),
    .O(\PCI-ROM/RC4 )
  );
  X_AND2   \PCI-ROM/$1I8219  (
    .I0(\PCI-ROM/SELA ),
    .I1(SUB_DATA5),
    .O(\PCI-ROM/RC5 )
  );
  X_AND2   \PCI-ROM/$1I8218  (
    .I0(\PCI-ROM/SELA ),
    .I1(SUB_DATA6),
    .O(\PCI-ROM/RC6 )
  );
  X_AND2   \PCI-ROM/$1I8217  (
    .I0(\PCI-ROM/SELA ),
    .I1(SUB_DATA7),
    .O(\PCI-ROM/RC7 )
  );
  X_AND2   \PCI-ROM/$1I8216  (
    .I0(\PCI-ROM/SELA ),
    .I1(SUB_DATA8),
    .O(\PCI-ROM/RC8 )
  );
  X_AND2   \PCI-ROM/$1I8215  (
    .I0(\PCI-ROM/SELA ),
    .I1(SUB_DATA9),
    .O(\PCI-ROM/RC9 )
  );
  X_AND2   \PCI-ROM/$1I8214  (
    .I0(\PCI-ROM/SELA ),
    .I1(SUB_DATA10),
    .O(\PCI-ROM/RC10 )
  );
  X_AND2   \PCI-ROM/$1I8213  (
    .I0(\PCI-ROM/SELA ),
    .I1(SUB_DATA11),
    .O(\PCI-ROM/RC11 )
  );
  X_AND2   \PCI-ROM/$1I8212  (
    .I0(\PCI-ROM/SELA ),
    .I1(SUB_DATA12),
    .O(\PCI-ROM/RC12 )
  );
  X_AND2   \PCI-ROM/$1I8211  (
    .I0(\PCI-ROM/SELA ),
    .I1(SUB_DATA13),
    .O(\PCI-ROM/RC13 )
  );
  X_AND2   \PCI-ROM/$1I8210  (
    .I0(\PCI-ROM/SELA ),
    .I1(SUB_DATA14),
    .O(\PCI-ROM/RC14 )
  );
  X_AND2   \PCI-ROM/$1I8209  (
    .I0(\PCI-ROM/SELA ),
    .I1(SUB_DATA15),
    .O(\PCI-ROM/RC15 )
  );
  X_AND2   \PCI-ROM/$1I8208  (
    .I0(\PCI-ROM/SELA ),
    .I1(SUB_DATA16),
    .O(\PCI-ROM/RC16 )
  );
  X_AND2   \PCI-ROM/$1I8207  (
    .I0(\PCI-ROM/SELA ),
    .I1(SUB_DATA17),
    .O(\PCI-ROM/RC17 )
  );
  X_AND2   \PCI-ROM/$1I8206  (
    .I0(\PCI-ROM/SELA ),
    .I1(SUB_DATA18),
    .O(\PCI-ROM/RC18 )
  );
  X_AND2   \PCI-ROM/$1I8205  (
    .I0(\PCI-ROM/SELA ),
    .I1(SUB_DATA19),
    .O(\PCI-ROM/RC19 )
  );
  X_AND2   \PCI-ROM/$1I8204  (
    .I0(\PCI-ROM/SELA ),
    .I1(SUB_DATA20),
    .O(\PCI-ROM/RC20 )
  );
  X_AND2   \PCI-ROM/$1I8203  (
    .I0(\PCI-ROM/SELA ),
    .I1(SUB_DATA21),
    .O(\PCI-ROM/RC21 )
  );
  X_AND2   \PCI-ROM/$1I8202  (
    .I0(\PCI-ROM/SELA ),
    .I1(SUB_DATA22),
    .O(\PCI-ROM/RC22 )
  );
  X_AND2   \PCI-ROM/$1I8201  (
    .I0(\PCI-ROM/SELA ),
    .I1(SUB_DATA23),
    .O(\PCI-ROM/RC23 )
  );
  X_AND2   \PCI-ROM/$1I8200  (
    .I0(\PCI-ROM/SELA ),
    .I1(SUB_DATA24),
    .O(\PCI-ROM/RC24 )
  );
  X_AND2   \PCI-ROM/$1I8199  (
    .I0(\PCI-ROM/SELA ),
    .I1(SUB_DATA25),
    .O(\PCI-ROM/RC25 )
  );
  X_AND2   \PCI-ROM/$1I8198  (
    .I0(\PCI-ROM/SELA ),
    .I1(SUB_DATA26),
    .O(\PCI-ROM/RC26 )
  );
  X_AND2   \PCI-ROM/$1I8197  (
    .I0(\PCI-ROM/SELA ),
    .I1(SUB_DATA27),
    .O(\PCI-ROM/RC27 )
  );
  X_AND2   \PCI-ROM/$1I8196  (
    .I0(\PCI-ROM/SELA ),
    .I1(SUB_DATA28),
    .O(\PCI-ROM/RC28 )
  );
  X_AND2   \PCI-ROM/$1I8195  (
    .I0(\PCI-ROM/SELA ),
    .I1(SUB_DATA29),
    .O(\PCI-ROM/RC29 )
  );
  X_AND2   \PCI-ROM/$1I8194  (
    .I0(\PCI-ROM/SELA ),
    .I1(SUB_DATA30),
    .O(\PCI-ROM/RC30 )
  );
  X_AND2   \PCI-ROM/$1I8193  (
    .I0(\PCI-ROM/SELA ),
    .I1(SUB_DATA31),
    .O(\PCI-ROM/RC31 )
  );
  X_AND2   \PCI-ROM/$1I8180  (
    .I0(\PCI-ROM/SEL0 ),
    .I1(CFG120),
    .O(\PCI-ROM/RA0 )
  );
  X_AND2   \PCI-ROM/$1I8179  (
    .I0(\PCI-ROM/SEL0 ),
    .I1(CFG121),
    .O(\PCI-ROM/RA1 )
  );
  X_AND2   \PCI-ROM/$1I8178  (
    .I0(\PCI-ROM/SEL0 ),
    .I1(CFG122),
    .O(\PCI-ROM/RA2 )
  );
  X_AND2   \PCI-ROM/$1I8177  (
    .I0(\PCI-ROM/SEL0 ),
    .I1(CFG123),
    .O(\PCI-ROM/RA3 )
  );
  X_AND2   \PCI-ROM/$1I8176  (
    .I0(\PCI-ROM/SEL0 ),
    .I1(CFG124),
    .O(\PCI-ROM/RA4 )
  );
  X_AND2   \PCI-ROM/$1I8175  (
    .I0(\PCI-ROM/SEL0 ),
    .I1(CFG125),
    .O(\PCI-ROM/RA5 )
  );
  X_AND2   \PCI-ROM/$1I8174  (
    .I0(\PCI-ROM/SEL0 ),
    .I1(CFG126),
    .O(\PCI-ROM/RA6 )
  );
  X_AND2   \PCI-ROM/$1I8173  (
    .I0(\PCI-ROM/SEL0 ),
    .I1(CFG127),
    .O(\PCI-ROM/RA7 )
  );
  X_AND2   \PCI-ROM/$1I8172  (
    .I0(\PCI-ROM/SEL0 ),
    .I1(CFG128),
    .O(\PCI-ROM/RA8 )
  );
  X_AND2   \PCI-ROM/$1I8171  (
    .I0(\PCI-ROM/SEL0 ),
    .I1(CFG129),
    .O(\PCI-ROM/RA9 )
  );
  X_AND2   \PCI-ROM/$1I8170  (
    .I0(\PCI-ROM/SEL0 ),
    .I1(CFG130),
    .O(\PCI-ROM/RA10 )
  );
  X_AND2   \PCI-ROM/$1I8169  (
    .I0(\PCI-ROM/SEL0 ),
    .I1(CFG131),
    .O(\PCI-ROM/RA11 )
  );
  X_AND2   \PCI-ROM/$1I8168  (
    .I0(\PCI-ROM/SEL0 ),
    .I1(CFG132),
    .O(\PCI-ROM/RA12 )
  );
  X_AND2   \PCI-ROM/$1I8167  (
    .I0(\PCI-ROM/SEL0 ),
    .I1(CFG133),
    .O(\PCI-ROM/RA13 )
  );
  X_AND2   \PCI-ROM/$1I8166  (
    .I0(\PCI-ROM/SEL0 ),
    .I1(CFG134),
    .O(\PCI-ROM/RA14 )
  );
  X_AND2   \PCI-ROM/$1I8165  (
    .I0(\PCI-ROM/SEL0 ),
    .I1(CFG135),
    .O(\PCI-ROM/RA15 )
  );
  X_AND2   \PCI-ROM/$1I8164  (
    .I0(\PCI-ROM/SEL0 ),
    .I1(CFG136),
    .O(\PCI-ROM/RA16 )
  );
  X_AND2   \PCI-ROM/$1I8163  (
    .I0(\PCI-ROM/SEL0 ),
    .I1(CFG137),
    .O(\PCI-ROM/RA17 )
  );
  X_AND2   \PCI-ROM/$1I8162  (
    .I0(\PCI-ROM/SEL0 ),
    .I1(CFG138),
    .O(\PCI-ROM/RA18 )
  );
  X_AND2   \PCI-ROM/$1I8161  (
    .I0(\PCI-ROM/SEL0 ),
    .I1(CFG139),
    .O(\PCI-ROM/RA19 )
  );
  X_AND2   \PCI-ROM/$1I8160  (
    .I0(\PCI-ROM/SEL0 ),
    .I1(CFG140),
    .O(\PCI-ROM/RA20 )
  );
  X_AND2   \PCI-ROM/$1I8159  (
    .I0(\PCI-ROM/SEL0 ),
    .I1(CFG141),
    .O(\PCI-ROM/RA21 )
  );
  X_AND2   \PCI-ROM/$1I8158  (
    .I0(\PCI-ROM/SEL0 ),
    .I1(CFG142),
    .O(\PCI-ROM/RA22 )
  );
  X_AND2   \PCI-ROM/$1I8157  (
    .I0(\PCI-ROM/SEL0 ),
    .I1(CFG143),
    .O(\PCI-ROM/RA23 )
  );
  X_AND2   \PCI-ROM/$1I8156  (
    .I0(\PCI-ROM/SEL0 ),
    .I1(CFG144),
    .O(\PCI-ROM/RA24 )
  );
  X_AND2   \PCI-ROM/$1I8155  (
    .I0(\PCI-ROM/SEL0 ),
    .I1(CFG145),
    .O(\PCI-ROM/RA25 )
  );
  X_AND2   \PCI-ROM/$1I8154  (
    .I0(\PCI-ROM/SEL0 ),
    .I1(CFG146),
    .O(\PCI-ROM/RA26 )
  );
  X_AND2   \PCI-ROM/$1I8153  (
    .I0(\PCI-ROM/SEL0 ),
    .I1(CFG147),
    .O(\PCI-ROM/RA27 )
  );
  X_AND2   \PCI-ROM/$1I8152  (
    .I0(\PCI-ROM/SEL0 ),
    .I1(CFG148),
    .O(\PCI-ROM/RA28 )
  );
  X_AND2   \PCI-ROM/$1I8151  (
    .I0(\PCI-ROM/SEL0 ),
    .I1(CFG149),
    .O(\PCI-ROM/RA29 )
  );
  X_AND2   \PCI-ROM/$1I8150  (
    .I0(\PCI-ROM/SEL0 ),
    .I1(CFG150),
    .O(\PCI-ROM/RA30 )
  );
  X_AND2   \PCI-ROM/$1I8149  (
    .I0(\PCI-ROM/SEL0 ),
    .I1(CFG151),
    .O(\PCI-ROM/RA31 )
  );
  X_AND2   \PCI-ROM/$1I8148  (
    .I0(\PCI-ROM/SEL2 ),
    .I1(CFG152),
    .O(\PCI-ROM/RB0 )
  );
  X_AND2   \PCI-ROM/$1I8147  (
    .I0(\PCI-ROM/SEL2 ),
    .I1(CFG153),
    .O(\PCI-ROM/RB1 )
  );
  X_AND2   \PCI-ROM/$1I8146  (
    .I0(\PCI-ROM/SEL2 ),
    .I1(CFG154),
    .O(\PCI-ROM/RB2 )
  );
  X_AND2   \PCI-ROM/$1I8145  (
    .I0(\PCI-ROM/SEL2 ),
    .I1(CFG155),
    .O(\PCI-ROM/RB3 )
  );
  X_AND2   \PCI-ROM/$1I8144  (
    .I0(\PCI-ROM/SEL2 ),
    .I1(CFG156),
    .O(\PCI-ROM/RB4 )
  );
  X_AND2   \PCI-ROM/$1I8143  (
    .I0(\PCI-ROM/SEL2 ),
    .I1(CFG157),
    .O(\PCI-ROM/RB5 )
  );
  X_AND2   \PCI-ROM/$1I8142  (
    .I0(\PCI-ROM/SEL2 ),
    .I1(CFG158),
    .O(\PCI-ROM/RB6 )
  );
  X_AND2   \PCI-ROM/$1I8141  (
    .I0(\PCI-ROM/SEL2 ),
    .I1(CFG159),
    .O(\PCI-ROM/RB7 )
  );
  X_AND2   \PCI-ROM/$1I8140  (
    .I0(\PCI-ROM/SEL2 ),
    .I1(CFG160),
    .O(\PCI-ROM/RB8 )
  );
  X_AND2   \PCI-ROM/$1I8139  (
    .I0(\PCI-ROM/SEL2 ),
    .I1(CFG161),
    .O(\PCI-ROM/RB9 )
  );
  X_AND2   \PCI-ROM/$1I8138  (
    .I0(\PCI-ROM/SEL2 ),
    .I1(CFG162),
    .O(\PCI-ROM/RB10 )
  );
  X_AND2   \PCI-ROM/$1I8137  (
    .I0(\PCI-ROM/SEL2 ),
    .I1(CFG163),
    .O(\PCI-ROM/RB11 )
  );
  X_AND2   \PCI-ROM/$1I8136  (
    .I0(\PCI-ROM/SEL2 ),
    .I1(CFG164),
    .O(\PCI-ROM/RB12 )
  );
  X_AND2   \PCI-ROM/$1I8135  (
    .I0(\PCI-ROM/SEL2 ),
    .I1(CFG165),
    .O(\PCI-ROM/RB13 )
  );
  X_AND2   \PCI-ROM/$1I8134  (
    .I0(\PCI-ROM/SEL2 ),
    .I1(CFG166),
    .O(\PCI-ROM/RB14 )
  );
  X_AND2   \PCI-ROM/$1I8133  (
    .I0(\PCI-ROM/SEL2 ),
    .I1(CFG167),
    .O(\PCI-ROM/RB15 )
  );
  X_AND2   \PCI-ROM/$1I8132  (
    .I0(\PCI-ROM/SEL2 ),
    .I1(CFG168),
    .O(\PCI-ROM/RB16 )
  );
  X_AND2   \PCI-ROM/$1I8131  (
    .I0(\PCI-ROM/SEL2 ),
    .I1(CFG169),
    .O(\PCI-ROM/RB17 )
  );
  X_AND2   \PCI-ROM/$1I8130  (
    .I0(\PCI-ROM/SEL2 ),
    .I1(CFG170),
    .O(\PCI-ROM/RB18 )
  );
  X_AND2   \PCI-ROM/$1I8129  (
    .I0(\PCI-ROM/SEL2 ),
    .I1(CFG171),
    .O(\PCI-ROM/RB19 )
  );
  X_AND2   \PCI-ROM/$1I8128  (
    .I0(\PCI-ROM/SEL2 ),
    .I1(CFG172),
    .O(\PCI-ROM/RB20 )
  );
  X_AND2   \PCI-ROM/$1I8127  (
    .I0(\PCI-ROM/SEL2 ),
    .I1(CFG173),
    .O(\PCI-ROM/RB21 )
  );
  X_AND2   \PCI-ROM/$1I8126  (
    .I0(\PCI-ROM/SEL2 ),
    .I1(CFG174),
    .O(\PCI-ROM/RB22 )
  );
  X_AND2   \PCI-ROM/$1I8125  (
    .I0(\PCI-ROM/SEL2 ),
    .I1(CFG175),
    .O(\PCI-ROM/RB23 )
  );
  X_AND2   \PCI-ROM/$1I8124  (
    .I0(\PCI-ROM/SEL2 ),
    .I1(CFG176),
    .O(\PCI-ROM/RB24 )
  );
  X_AND2   \PCI-ROM/$1I8123  (
    .I0(\PCI-ROM/SEL2 ),
    .I1(CFG177),
    .O(\PCI-ROM/RB25 )
  );
  X_AND2   \PCI-ROM/$1I8122  (
    .I0(\PCI-ROM/SEL2 ),
    .I1(CFG178),
    .O(\PCI-ROM/RB26 )
  );
  X_AND2   \PCI-ROM/$1I8121  (
    .I0(\PCI-ROM/SEL2 ),
    .I1(CFG179),
    .O(\PCI-ROM/RB27 )
  );
  X_AND2   \PCI-ROM/$1I8120  (
    .I0(\PCI-ROM/SEL2 ),
    .I1(CFG180),
    .O(\PCI-ROM/RB28 )
  );
  X_AND2   \PCI-ROM/$1I8119  (
    .I0(\PCI-ROM/SEL2 ),
    .I1(CFG181),
    .O(\PCI-ROM/RB29 )
  );
  X_AND2   \PCI-ROM/$1I8118  (
    .I0(\PCI-ROM/SEL2 ),
    .I1(CFG182),
    .O(\PCI-ROM/RB30 )
  );
  X_AND2   \PCI-ROM/$1I8117  (
    .I0(\PCI-ROM/SEL2 ),
    .I1(CFG183),
    .O(\PCI-ROM/RB31 )
  );
  X_AND3   \PCI-ROM/$1I8110  (
    .I0(\NlwInverterSignal_PCI-ROM/$1I8110/I0 ),
    .I1(\NlwInverterSignal_PCI-ROM/$1I8110/I1 ),
    .I2(\PCI-ROM/$1N8111 ),
    .O(\PCI-ROM/SEL2 )
  );
  X_AND3   \PCI-ROM/$1I8078  (
    .I0(\NlwInverterSignal_PCI-ROM/$1I8078/I0 ),
    .I1(\NlwInverterSignal_PCI-ROM/$1I8078/I1 ),
    .I2(\PCI-ROM/$1N7806 ),
    .O(\PCI-ROM/SEL0 )
  );
  X_AND4   \PCI-ROM/$1I7800/AND4  (
    .I0(\PCI-ROM/$1I7800/$1N2275 ),
    .I1(\PCI-ROM/$1I7800/$1N2276 ),
    .I2(\PCI-ROM/$1I7800/$1N2277 ),
    .I3(\PCI-ROM/$1I7800/$1N2283 ),
    .O(\PCI-ROM/$1N7806 )
  );
  X_INV   \PCI-ROM/$1I7800/INV3  (
    .I(NlwRenamedSig_OI_ADDR5),
    .O(\PCI-ROM/$1I7800/$1N2283 )
  );
  X_INV   \PCI-ROM/$1I7800/INV2  (
    .I(NlwRenamedSig_OI_ADDR4),
    .O(\PCI-ROM/$1I7800/$1N2277 )
  );
  X_INV   \PCI-ROM/$1I7800/INV1  (
    .I(NlwRenamedSig_OI_ADDR3),
    .O(\PCI-ROM/$1I7800/$1N2276 )
  );
  X_INV   \PCI-ROM/$1I7800/INV0  (
    .I(NlwRenamedSig_OI_ADDR2),
    .O(\PCI-ROM/$1I7800/$1N2275 )
  );
  X_AND4   \PCI-ROM/$1I8181/AND4  (
    .I0(\PCI-ROM/$1I8181/$1N2275 ),
    .I1(NlwRenamedSig_OI_ADDR3),
    .I2(\PCI-ROM/$1I8181/$1N2277 ),
    .I3(\PCI-ROM/$1I8181/$1N2283 ),
    .O(\PCI-ROM/$1N8111 )
  );
  X_INV   \PCI-ROM/$1I8181/INV3  (
    .I(NlwRenamedSig_OI_ADDR5),
    .O(\PCI-ROM/$1I8181/$1N2283 )
  );
  X_INV   \PCI-ROM/$1I8181/INV2  (
    .I(NlwRenamedSig_OI_ADDR4),
    .O(\PCI-ROM/$1I8181/$1N2277 )
  );
  X_INV   \PCI-ROM/$1I8181/INV0  (
    .I(NlwRenamedSig_OI_ADDR2),
    .O(\PCI-ROM/$1I8181/$1N2275 )
  );
  X_AND4   \PCI-ROM/$1I8225/AND4  (
    .I0(\PCI-ROM/$1I8225/$1N2275 ),
    .I1(NlwRenamedSig_OI_ADDR3),
    .I2(\PCI-ROM/$1I8225/$1N2277 ),
    .I3(NlwRenamedSig_OI_ADDR5),
    .O(\PCI-ROM/$1N8188 )
  );
  X_INV   \PCI-ROM/$1I8225/INV2  (
    .I(NlwRenamedSig_OI_ADDR4),
    .O(\PCI-ROM/$1I8225/$1N2277 )
  );
  X_INV   \PCI-ROM/$1I8225/INV0  (
    .I(NlwRenamedSig_OI_ADDR2),
    .O(\PCI-ROM/$1I8225/$1N2275 )
  );
  X_AND4   \PCI-ROM/$1I8276/AND4  (
    .I0(NlwRenamedSig_OI_ADDR2),
    .I1(NlwRenamedSig_OI_ADDR3),
    .I2(\PCI-ROM/$1I8276/$1N2277 ),
    .I3(NlwRenamedSig_OI_ADDR5),
    .O(\PCI-ROM/$1N8238 )
  );
  X_INV   \PCI-ROM/$1I8276/INV2  (
    .I(NlwRenamedSig_OI_ADDR4),
    .O(\PCI-ROM/$1I8276/$1N2277 )
  );
  X_AND4   \PCI-ROM/$1I8288/AND4  (
    .I0(NlwRenamedSig_OI_ADDR2),
    .I1(NlwRenamedSig_OI_ADDR3),
    .I2(\PCI-ROM/$1I8288/$1N2277 ),
    .I3(NlwRenamedSig_OI_ADDR5),
    .O(\PCI-ROM/$1N8283 )
  );
  X_INV   \PCI-ROM/$1I8288/INV2  (
    .I(NlwRenamedSig_OI_ADDR4),
    .O(\PCI-ROM/$1I8288/$1N2277 )
  );
  X_AND4   \PCI-ROM/$1I8332/AND4  (
    .I0(NlwRenamedSig_OI_ADDR2),
    .I1(\PCI-ROM/$1I8332/$1N2290 ),
    .I2(NlwRenamedSig_OI_ADDR4),
    .I3(NlwRenamedSig_OI_ADDR5),
    .O(\PCI-ROM/$1N8328 )
  );
  X_INV   \PCI-ROM/$1I8332/INV1  (
    .I(NlwRenamedSig_OI_ADDR3),
    .O(\PCI-ROM/$1I8332/$1N2290 )
  );
  X_ZERO   \PCI-ROM/$1I8452/$1I2218  (
    .O(\PCI-ROM/$1I8452/$1N2216 )
  );
  X_BUF   \PCI-ROM/$1I8452/L  (
    .I(\PCI-ROM/$1I8452/$1N2216 ),
    .O(\PCI-ROM/$1N8453 )
  );
  X_BUF   \PCI-ROM/$1I8479/NC  (
    .I(\PCI-ROM/CLR31 ),
    .O(\NLW_PCI-ROM/$1I8479/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-ROM/$1I8480/NC  (
    .I(\PCI-ROM/CLR30 ),
    .O(\NLW_PCI-ROM/$1I8480/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-ROM/$1I8481/NC  (
    .I(\PCI-ROM/CLR29 ),
    .O(\NLW_PCI-ROM/$1I8481/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-ROM/$1I8482/NC  (
    .I(\PCI-ROM/CLR28 ),
    .O(\NLW_PCI-ROM/$1I8482/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-ROM/$1I8483/NC  (
    .I(\PCI-ROM/CLR27 ),
    .O(\NLW_PCI-ROM/$1I8483/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-ROM/$1I8484/NC  (
    .I(\PCI-ROM/CLR26 ),
    .O(\NLW_PCI-ROM/$1I8484/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-ROM/$1I8485/NC  (
    .I(\PCI-ROM/CLR25 ),
    .O(\NLW_PCI-ROM/$1I8485/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-ROM/$1I8486/NC  (
    .I(\PCI-ROM/CLR24 ),
    .O(\NLW_PCI-ROM/$1I8486/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-ROM/$1I8487/NC  (
    .I(\PCI-ROM/CLR23 ),
    .O(\NLW_PCI-ROM/$1I8487/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-ROM/$1I8488/NC  (
    .I(\PCI-ROM/CLR22 ),
    .O(\NLW_PCI-ROM/$1I8488/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-ROM/$1I8489/NC  (
    .I(\PCI-ROM/CLR21 ),
    .O(\NLW_PCI-ROM/$1I8489/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-ROM/$1I8490/NC  (
    .I(\PCI-ROM/CLR20 ),
    .O(\NLW_PCI-ROM/$1I8490/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-ROM/$1I8491/NC  (
    .I(\PCI-ROM/CLR19 ),
    .O(\NLW_PCI-ROM/$1I8491/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-ROM/$1I8492/NC  (
    .I(\PCI-ROM/CLR18 ),
    .O(\NLW_PCI-ROM/$1I8492/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-ROM/$1I8493/NC  (
    .I(\PCI-ROM/CLR17 ),
    .O(\NLW_PCI-ROM/$1I8493/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-ROM/$1I8494/NC  (
    .I(\PCI-ROM/CLR16 ),
    .O(\NLW_PCI-ROM/$1I8494/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-ROM/$1I8495/NC  (
    .I(\PCI-ROM/CLR15 ),
    .O(\NLW_PCI-ROM/$1I8495/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-ROM/$1I8496/NC  (
    .I(\PCI-ROM/CLR14 ),
    .O(\NLW_PCI-ROM/$1I8496/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-ROM/$1I8497/NC  (
    .I(\PCI-ROM/CLR13 ),
    .O(\NLW_PCI-ROM/$1I8497/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-ROM/$1I8498/NC  (
    .I(\PCI-ROM/CLR12 ),
    .O(\NLW_PCI-ROM/$1I8498/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-ROM/$1I8499/NC  (
    .I(\PCI-ROM/CLR11 ),
    .O(\NLW_PCI-ROM/$1I8499/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-ROM/$1I8500/NC  (
    .I(\PCI-ROM/CLR10 ),
    .O(\NLW_PCI-ROM/$1I8500/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-ROM/$1I8501/NC  (
    .I(\PCI-ROM/CLR9 ),
    .O(\NLW_PCI-ROM/$1I8501/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-ROM/$1I8502/NC  (
    .I(\PCI-ROM/CLR8 ),
    .O(\NLW_PCI-ROM/$1I8502/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-ROM/$1I8503/NC  (
    .I(\PCI-ROM/CLR7 ),
    .O(\NLW_PCI-ROM/$1I8503/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-ROM/$1I8504/NC  (
    .I(\PCI-ROM/CLR6 ),
    .O(\NLW_PCI-ROM/$1I8504/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-ROM/$1I8505/NC  (
    .I(\PCI-ROM/CLR5 ),
    .O(\NLW_PCI-ROM/$1I8505/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-ROM/$1I8506/NC  (
    .I(\PCI-ROM/CLR4 ),
    .O(\NLW_PCI-ROM/$1I8506/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-ROM/$1I8507/NC  (
    .I(\PCI-ROM/CLR3 ),
    .O(\NLW_PCI-ROM/$1I8507/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-ROM/$1I8508/NC  (
    .I(\PCI-ROM/CLR2 ),
    .O(\NLW_PCI-ROM/$1I8508/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-ROM/$1I8509/NC  (
    .I(\PCI-ROM/CLR1 ),
    .O(\NLW_PCI-ROM/$1I8509/NC_O_UNCONNECTED )
  );
  X_BUF   \PCI-ROM/$1I8510/NC  (
    .I(\PCI-ROM/CLR0 ),
    .O(\NLW_PCI-ROM/$1I8510/NC_O_UNCONNECTED )
  );
  X_INV   \$4I4029/$1I2779  (
    .I(\$4I4029/ONE ),
    .O(\$4I4029/$1N2778 )
  );
  X_AND2   \$4I4029/$1I2776  (
    .I0(\$4I4029/$1N2763 ),
    .I1(\$4I4029/$1N2778 ),
    .O(EX)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \$4I4029/$1I2756  (
    .CLK(CLK),
    .I(\$4I4029/$1N2757 ),
    .O(\$4I4029/$1N2759 ),
    .RST(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \$4I4029/$1I2752  (
    .CLK(CLK),
    .I(\$4I4029/$1N2753 ),
    .O(\$4I4029/$1N2755 ),
    .RST(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \$4I4029/$1I2748  (
    .CLK(CLK),
    .I(\$4I4029/$1N2749 ),
    .O(\$4I4029/$1N2751 ),
    .RST(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \$4I4029/$1I2732  (
    .CLK(CLK),
    .I(\$4I4029/$1N2711 ),
    .O(\$4I4029/$1N2734 ),
    .RST(NlwRenamedSig_OI_RST),
    .CE(VCC),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \$4I4029/$1I2725  (
    .CE(\$4I4029/EXP ),
    .CLK(CLK),
    .I(\$4I4029/ONE ),
    .O(\$4I4029/$1N2763 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND2   \$4I4029/$1I2610/$1I31  (
    .I0(\$4I4029/$1N2616 ),
    .I1(\$4I4029/$1I2610/TC ),
    .O(\$4I4029/$1N2711 )
  );
  X_AND4   \$4I4029/$1I2610/$1I28  (
    .I0(\$4I4029/$1I2610/Q6 ),
    .I1(\$4I4029/$1I2610/Q5 ),
    .I2(\$4I4029/$1I2610/Q4 ),
    .I3(\$4I4029/$1I2610/T4 ),
    .O(\$4I4029/$1I2610/T7 )
  );
  X_AND3   \$4I4029/$1I2610/$1I26  (
    .I0(\$4I4029/$1I2610/Q2 ),
    .I1(\$4I4029/$1I2610/Q1 ),
    .I2(\$4I4029/$1I2610/Q0 ),
    .O(\$4I4029/$1I2610/T3 )
  );
  X_AND2   \$4I4029/$1I2610/$1I24  (
    .I0(\$4I4029/$1I2610/Q1 ),
    .I1(\$4I4029/$1I2610/Q0 ),
    .O(\$4I4029/$1I2610/T2 )
  );
  X_AND2   \$4I4029/$1I2610/$1I2  (
    .I0(\$4I4029/$1I2610/Q4 ),
    .I1(\$4I4029/$1I2610/T4 ),
    .O(\$4I4029/$1I2610/T5 )
  );
  X_ONE   \$4I4029/$1I2610/$1I16  (
    .O(\$4I4029/$1I2610/$1N20 )
  );
  X_AND4   \$4I4029/$1I2610/$1I15  (
    .I0(\$4I4029/$1I2610/Q3 ),
    .I1(\$4I4029/$1I2610/Q2 ),
    .I2(\$4I4029/$1I2610/Q1 ),
    .I3(\$4I4029/$1I2610/Q0 ),
    .O(\$4I4029/$1I2610/T4 )
  );
  X_AND3   \$4I4029/$1I2610/$1I11  (
    .I0(\$4I4029/$1I2610/Q5 ),
    .I1(\$4I4029/$1I2610/Q4 ),
    .I2(\$4I4029/$1I2610/T4 ),
    .O(\$4I4029/$1I2610/T6 )
  );
  X_AND5   \$4I4029/$1I2610/$1I1  (
    .I0(\$4I4029/$1I2610/Q7 ),
    .I1(\$4I4029/$1I2610/Q6 ),
    .I2(\$4I4029/$1I2610/Q5 ),
    .I3(\$4I4029/$1I2610/Q4 ),
    .I4(\$4I4029/$1I2610/T4 ),
    .O(\$4I4029/$1I2610/TC )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \$4I4029/$1I2610/$1I43/$1I35  (
    .CE(\$4I4029/$1N2616 ),
    .CLK(CLK),
    .I(\$4I4029/$1I2610/$1I43/MD ),
    .O(\$4I4029/$1I2610/Q0 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \$4I4029/$1I2610/$1I43/$1I32  (
    .I0(\$4I4029/$1I2610/$1N20 ),
    .I1(\$4I4029/$1I2610/Q0 ),
    .O(\$4I4029/$1I2610/$1I43/TQ )
  );
  X_AND2   \$4I4029/$1I2610/$1I43/$1I30/$1I9  (
    .I0(\$4I4029/$1I2610/$1N45 ),
    .I1(\$4I4029/$1I2610/$1N48 ),
    .O(\$4I4029/$1I2610/$1I43/$1I30/M1 )
  );
  X_OR2   \$4I4029/$1I2610/$1I43/$1I30/$1I8  (
    .I0(\$4I4029/$1I2610/$1I43/$1I30/M1 ),
    .I1(\$4I4029/$1I2610/$1I43/$1I30/M0 ),
    .O(\$4I4029/$1I2610/$1I43/MD )
  );
  X_AND2   \$4I4029/$1I2610/$1I43/$1I30/$1I7  (
    .I0(\NlwInverterSignal_$4I4029/$1I2610/$1I43/$1I30/$1I7/I0 ),
    .I1(\$4I4029/$1I2610/$1I43/TQ ),
    .O(\$4I4029/$1I2610/$1I43/$1I30/M0 )
  );
  X_ZERO   \$4I4029/$1I2610/$1I44/$1I2218  (
    .O(\$4I4029/$1I2610/$1I44/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2610/$1I44/L  (
    .I(\$4I4029/$1I2610/$1I44/$1N2216 ),
    .O(\$4I4029/$1I2610/$1N45 )
  );
  X_ZERO   \$4I4029/$1I2610/$1I47/$1I2218  (
    .O(\$4I4029/$1I2610/$1I47/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2610/$1I47/L  (
    .I(\$4I4029/$1I2610/$1I47/$1N2216 ),
    .O(\$4I4029/$1I2610/$1N48 )
  );
  X_ZERO   \$4I4029/$1I2610/$1I49/$1I2218  (
    .O(\$4I4029/$1I2610/$1I49/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2610/$1I49/L  (
    .I(\$4I4029/$1I2610/$1I49/$1N2216 ),
    .O(\$4I4029/$1I2610/$1N50 )
  );
  X_ZERO   \$4I4029/$1I2610/$1I52/$1I2218  (
    .O(\$4I4029/$1I2610/$1I52/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2610/$1I52/L  (
    .I(\$4I4029/$1I2610/$1I52/$1N2216 ),
    .O(\$4I4029/$1I2610/$1N51 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \$4I4029/$1I2610/$1I53/$1I35  (
    .CE(\$4I4029/$1N2616 ),
    .CLK(CLK),
    .I(\$4I4029/$1I2610/$1I53/MD ),
    .O(\$4I4029/$1I2610/Q1 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \$4I4029/$1I2610/$1I53/$1I32  (
    .I0(\$4I4029/$1I2610/Q0 ),
    .I1(\$4I4029/$1I2610/Q1 ),
    .O(\$4I4029/$1I2610/$1I53/TQ )
  );
  X_AND2   \$4I4029/$1I2610/$1I53/$1I30/$1I9  (
    .I0(\$4I4029/$1I2610/$1N50 ),
    .I1(\$4I4029/$1I2610/$1N51 ),
    .O(\$4I4029/$1I2610/$1I53/$1I30/M1 )
  );
  X_OR2   \$4I4029/$1I2610/$1I53/$1I30/$1I8  (
    .I0(\$4I4029/$1I2610/$1I53/$1I30/M1 ),
    .I1(\$4I4029/$1I2610/$1I53/$1I30/M0 ),
    .O(\$4I4029/$1I2610/$1I53/MD )
  );
  X_AND2   \$4I4029/$1I2610/$1I53/$1I30/$1I7  (
    .I0(\NlwInverterSignal_$4I4029/$1I2610/$1I53/$1I30/$1I7/I0 ),
    .I1(\$4I4029/$1I2610/$1I53/TQ ),
    .O(\$4I4029/$1I2610/$1I53/$1I30/M0 )
  );
  X_ZERO   \$4I4029/$1I2610/$1I54/$1I2218  (
    .O(\$4I4029/$1I2610/$1I54/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2610/$1I54/L  (
    .I(\$4I4029/$1I2610/$1I54/$1N2216 ),
    .O(\$4I4029/$1I2610/$1N55 )
  );
  X_ZERO   \$4I4029/$1I2610/$1I57/$1I2218  (
    .O(\$4I4029/$1I2610/$1I57/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2610/$1I57/L  (
    .I(\$4I4029/$1I2610/$1I57/$1N2216 ),
    .O(\$4I4029/$1I2610/$1N56 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \$4I4029/$1I2610/$1I58/$1I35  (
    .CE(\$4I4029/$1N2616 ),
    .CLK(CLK),
    .I(\$4I4029/$1I2610/$1I58/MD ),
    .O(\$4I4029/$1I2610/Q2 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \$4I4029/$1I2610/$1I58/$1I32  (
    .I0(\$4I4029/$1I2610/T2 ),
    .I1(\$4I4029/$1I2610/Q2 ),
    .O(\$4I4029/$1I2610/$1I58/TQ )
  );
  X_AND2   \$4I4029/$1I2610/$1I58/$1I30/$1I9  (
    .I0(\$4I4029/$1I2610/$1N55 ),
    .I1(\$4I4029/$1I2610/$1N56 ),
    .O(\$4I4029/$1I2610/$1I58/$1I30/M1 )
  );
  X_OR2   \$4I4029/$1I2610/$1I58/$1I30/$1I8  (
    .I0(\$4I4029/$1I2610/$1I58/$1I30/M1 ),
    .I1(\$4I4029/$1I2610/$1I58/$1I30/M0 ),
    .O(\$4I4029/$1I2610/$1I58/MD )
  );
  X_AND2   \$4I4029/$1I2610/$1I58/$1I30/$1I7  (
    .I0(\NlwInverterSignal_$4I4029/$1I2610/$1I58/$1I30/$1I7/I0 ),
    .I1(\$4I4029/$1I2610/$1I58/TQ ),
    .O(\$4I4029/$1I2610/$1I58/$1I30/M0 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \$4I4029/$1I2610/$1I59/$1I35  (
    .CE(\$4I4029/$1N2616 ),
    .CLK(CLK),
    .I(\$4I4029/$1I2610/$1I59/MD ),
    .O(\$4I4029/$1I2610/Q3 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \$4I4029/$1I2610/$1I59/$1I32  (
    .I0(\$4I4029/$1I2610/T3 ),
    .I1(\$4I4029/$1I2610/Q3 ),
    .O(\$4I4029/$1I2610/$1I59/TQ )
  );
  X_AND2   \$4I4029/$1I2610/$1I59/$1I30/$1I9  (
    .I0(\$4I4029/$1I2610/$1N62 ),
    .I1(\$4I4029/$1I2610/$1N61 ),
    .O(\$4I4029/$1I2610/$1I59/$1I30/M1 )
  );
  X_OR2   \$4I4029/$1I2610/$1I59/$1I30/$1I8  (
    .I0(\$4I4029/$1I2610/$1I59/$1I30/M1 ),
    .I1(\$4I4029/$1I2610/$1I59/$1I30/M0 ),
    .O(\$4I4029/$1I2610/$1I59/MD )
  );
  X_AND2   \$4I4029/$1I2610/$1I59/$1I30/$1I7  (
    .I0(\NlwInverterSignal_$4I4029/$1I2610/$1I59/$1I30/$1I7/I0 ),
    .I1(\$4I4029/$1I2610/$1I59/TQ ),
    .O(\$4I4029/$1I2610/$1I59/$1I30/M0 )
  );
  X_ZERO   \$4I4029/$1I2610/$1I60/$1I2218  (
    .O(\$4I4029/$1I2610/$1I60/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2610/$1I60/L  (
    .I(\$4I4029/$1I2610/$1I60/$1N2216 ),
    .O(\$4I4029/$1I2610/$1N61 )
  );
  X_ZERO   \$4I4029/$1I2610/$1I63/$1I2218  (
    .O(\$4I4029/$1I2610/$1I63/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2610/$1I63/L  (
    .I(\$4I4029/$1I2610/$1I63/$1N2216 ),
    .O(\$4I4029/$1I2610/$1N62 )
  );
  X_ZERO   \$4I4029/$1I2610/$1I64/$1I2218  (
    .O(\$4I4029/$1I2610/$1I64/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2610/$1I64/L  (
    .I(\$4I4029/$1I2610/$1I64/$1N2216 ),
    .O(\$4I4029/$1I2610/$1N65 )
  );
  X_ZERO   \$4I4029/$1I2610/$1I67/$1I2218  (
    .O(\$4I4029/$1I2610/$1I67/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2610/$1I67/L  (
    .I(\$4I4029/$1I2610/$1I67/$1N2216 ),
    .O(\$4I4029/$1I2610/$1N66 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \$4I4029/$1I2610/$1I68/$1I35  (
    .CE(\$4I4029/$1N2616 ),
    .CLK(CLK),
    .I(\$4I4029/$1I2610/$1I68/MD ),
    .O(\$4I4029/$1I2610/Q4 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \$4I4029/$1I2610/$1I68/$1I32  (
    .I0(\$4I4029/$1I2610/T4 ),
    .I1(\$4I4029/$1I2610/Q4 ),
    .O(\$4I4029/$1I2610/$1I68/TQ )
  );
  X_AND2   \$4I4029/$1I2610/$1I68/$1I30/$1I9  (
    .I0(\$4I4029/$1I2610/$1N65 ),
    .I1(\$4I4029/$1I2610/$1N66 ),
    .O(\$4I4029/$1I2610/$1I68/$1I30/M1 )
  );
  X_OR2   \$4I4029/$1I2610/$1I68/$1I30/$1I8  (
    .I0(\$4I4029/$1I2610/$1I68/$1I30/M1 ),
    .I1(\$4I4029/$1I2610/$1I68/$1I30/M0 ),
    .O(\$4I4029/$1I2610/$1I68/MD )
  );
  X_AND2   \$4I4029/$1I2610/$1I68/$1I30/$1I7  (
    .I0(\NlwInverterSignal_$4I4029/$1I2610/$1I68/$1I30/$1I7/I0 ),
    .I1(\$4I4029/$1I2610/$1I68/TQ ),
    .O(\$4I4029/$1I2610/$1I68/$1I30/M0 )
  );
  X_ZERO   \$4I4029/$1I2610/$1I69/$1I2218  (
    .O(\$4I4029/$1I2610/$1I69/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2610/$1I69/L  (
    .I(\$4I4029/$1I2610/$1I69/$1N2216 ),
    .O(\$4I4029/$1I2610/$1N70 )
  );
  X_ZERO   \$4I4029/$1I2610/$1I72/$1I2218  (
    .O(\$4I4029/$1I2610/$1I72/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2610/$1I72/L  (
    .I(\$4I4029/$1I2610/$1I72/$1N2216 ),
    .O(\$4I4029/$1I2610/$1N71 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \$4I4029/$1I2610/$1I73/$1I35  (
    .CE(\$4I4029/$1N2616 ),
    .CLK(CLK),
    .I(\$4I4029/$1I2610/$1I73/MD ),
    .O(\$4I4029/$1I2610/Q5 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \$4I4029/$1I2610/$1I73/$1I32  (
    .I0(\$4I4029/$1I2610/T5 ),
    .I1(\$4I4029/$1I2610/Q5 ),
    .O(\$4I4029/$1I2610/$1I73/TQ )
  );
  X_AND2   \$4I4029/$1I2610/$1I73/$1I30/$1I9  (
    .I0(\$4I4029/$1I2610/$1N70 ),
    .I1(\$4I4029/$1I2610/$1N71 ),
    .O(\$4I4029/$1I2610/$1I73/$1I30/M1 )
  );
  X_OR2   \$4I4029/$1I2610/$1I73/$1I30/$1I8  (
    .I0(\$4I4029/$1I2610/$1I73/$1I30/M1 ),
    .I1(\$4I4029/$1I2610/$1I73/$1I30/M0 ),
    .O(\$4I4029/$1I2610/$1I73/MD )
  );
  X_AND2   \$4I4029/$1I2610/$1I73/$1I30/$1I7  (
    .I0(\NlwInverterSignal_$4I4029/$1I2610/$1I73/$1I30/$1I7/I0 ),
    .I1(\$4I4029/$1I2610/$1I73/TQ ),
    .O(\$4I4029/$1I2610/$1I73/$1I30/M0 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \$4I4029/$1I2610/$1I79/$1I35  (
    .CE(\$4I4029/$1N2616 ),
    .CLK(CLK),
    .I(\$4I4029/$1I2610/$1I79/MD ),
    .O(\$4I4029/$1I2610/Q6 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \$4I4029/$1I2610/$1I79/$1I32  (
    .I0(\$4I4029/$1I2610/T6 ),
    .I1(\$4I4029/$1I2610/Q6 ),
    .O(\$4I4029/$1I2610/$1I79/TQ )
  );
  X_AND2   \$4I4029/$1I2610/$1I79/$1I30/$1I9  (
    .I0(\$4I4029/$1I2610/$1N82 ),
    .I1(\$4I4029/$1I2610/$1N81 ),
    .O(\$4I4029/$1I2610/$1I79/$1I30/M1 )
  );
  X_OR2   \$4I4029/$1I2610/$1I79/$1I30/$1I8  (
    .I0(\$4I4029/$1I2610/$1I79/$1I30/M1 ),
    .I1(\$4I4029/$1I2610/$1I79/$1I30/M0 ),
    .O(\$4I4029/$1I2610/$1I79/MD )
  );
  X_AND2   \$4I4029/$1I2610/$1I79/$1I30/$1I7  (
    .I0(\NlwInverterSignal_$4I4029/$1I2610/$1I79/$1I30/$1I7/I0 ),
    .I1(\$4I4029/$1I2610/$1I79/TQ ),
    .O(\$4I4029/$1I2610/$1I79/$1I30/M0 )
  );
  X_ZERO   \$4I4029/$1I2610/$1I80/$1I2218  (
    .O(\$4I4029/$1I2610/$1I80/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2610/$1I80/L  (
    .I(\$4I4029/$1I2610/$1I80/$1N2216 ),
    .O(\$4I4029/$1I2610/$1N81 )
  );
  X_ZERO   \$4I4029/$1I2610/$1I83/$1I2218  (
    .O(\$4I4029/$1I2610/$1I83/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2610/$1I83/L  (
    .I(\$4I4029/$1I2610/$1I83/$1N2216 ),
    .O(\$4I4029/$1I2610/$1N82 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \$4I4029/$1I2610/$1I84/$1I35  (
    .CE(\$4I4029/$1N2616 ),
    .CLK(CLK),
    .I(\$4I4029/$1I2610/$1I84/MD ),
    .O(\$4I4029/$1I2610/Q7 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \$4I4029/$1I2610/$1I84/$1I32  (
    .I0(\$4I4029/$1I2610/T7 ),
    .I1(\$4I4029/$1I2610/Q7 ),
    .O(\$4I4029/$1I2610/$1I84/TQ )
  );
  X_AND2   \$4I4029/$1I2610/$1I84/$1I30/$1I9  (
    .I0(\$4I4029/$1I2610/$1N87 ),
    .I1(\$4I4029/$1I2610/$1N86 ),
    .O(\$4I4029/$1I2610/$1I84/$1I30/M1 )
  );
  X_OR2   \$4I4029/$1I2610/$1I84/$1I30/$1I8  (
    .I0(\$4I4029/$1I2610/$1I84/$1I30/M1 ),
    .I1(\$4I4029/$1I2610/$1I84/$1I30/M0 ),
    .O(\$4I4029/$1I2610/$1I84/MD )
  );
  X_AND2   \$4I4029/$1I2610/$1I84/$1I30/$1I7  (
    .I0(\NlwInverterSignal_$4I4029/$1I2610/$1I84/$1I30/$1I7/I0 ),
    .I1(\$4I4029/$1I2610/$1I84/TQ ),
    .O(\$4I4029/$1I2610/$1I84/$1I30/M0 )
  );
  X_ZERO   \$4I4029/$1I2610/$1I85/$1I2218  (
    .O(\$4I4029/$1I2610/$1I85/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2610/$1I85/L  (
    .I(\$4I4029/$1I2610/$1I85/$1N2216 ),
    .O(\$4I4029/$1I2610/$1N86 )
  );
  X_ZERO   \$4I4029/$1I2610/$1I88/$1I2218  (
    .O(\$4I4029/$1I2610/$1I88/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2610/$1I88/L  (
    .I(\$4I4029/$1I2610/$1I88/$1N2216 ),
    .O(\$4I4029/$1I2610/$1N87 )
  );
  X_ONE   \$4I4029/$1I2615/$1I2220  (
    .O(\$4I4029/$1I2615/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2615/H  (
    .I(\$4I4029/$1I2615/$1N2216 ),
    .O(\$4I4029/$1N2616 )
  );
  X_AND2   \$4I4029/$1I2637/$1I31  (
    .I0(\$4I4029/$1N2734 ),
    .I1(\$4I4029/$1I2637/TC ),
    .O(\$4I4029/$1N2749 )
  );
  X_AND4   \$4I4029/$1I2637/$1I28  (
    .I0(\$4I4029/$1I2637/Q6 ),
    .I1(\$4I4029/$1I2637/Q5 ),
    .I2(\$4I4029/$1I2637/Q4 ),
    .I3(\$4I4029/$1I2637/T4 ),
    .O(\$4I4029/$1I2637/T7 )
  );
  X_AND3   \$4I4029/$1I2637/$1I26  (
    .I0(\$4I4029/$1I2637/Q2 ),
    .I1(\$4I4029/$1I2637/Q1 ),
    .I2(\$4I4029/$1I2637/Q0 ),
    .O(\$4I4029/$1I2637/T3 )
  );
  X_AND2   \$4I4029/$1I2637/$1I24  (
    .I0(\$4I4029/$1I2637/Q1 ),
    .I1(\$4I4029/$1I2637/Q0 ),
    .O(\$4I4029/$1I2637/T2 )
  );
  X_AND2   \$4I4029/$1I2637/$1I2  (
    .I0(\$4I4029/$1I2637/Q4 ),
    .I1(\$4I4029/$1I2637/T4 ),
    .O(\$4I4029/$1I2637/T5 )
  );
  X_ONE   \$4I4029/$1I2637/$1I16  (
    .O(\$4I4029/$1I2637/$1N20 )
  );
  X_AND4   \$4I4029/$1I2637/$1I15  (
    .I0(\$4I4029/$1I2637/Q3 ),
    .I1(\$4I4029/$1I2637/Q2 ),
    .I2(\$4I4029/$1I2637/Q1 ),
    .I3(\$4I4029/$1I2637/Q0 ),
    .O(\$4I4029/$1I2637/T4 )
  );
  X_AND3   \$4I4029/$1I2637/$1I11  (
    .I0(\$4I4029/$1I2637/Q5 ),
    .I1(\$4I4029/$1I2637/Q4 ),
    .I2(\$4I4029/$1I2637/T4 ),
    .O(\$4I4029/$1I2637/T6 )
  );
  X_AND5   \$4I4029/$1I2637/$1I1  (
    .I0(\$4I4029/$1I2637/Q7 ),
    .I1(\$4I4029/$1I2637/Q6 ),
    .I2(\$4I4029/$1I2637/Q5 ),
    .I3(\$4I4029/$1I2637/Q4 ),
    .I4(\$4I4029/$1I2637/T4 ),
    .O(\$4I4029/$1I2637/TC )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \$4I4029/$1I2637/$1I43/$1I35  (
    .CE(\$4I4029/$1N2734 ),
    .CLK(CLK),
    .I(\$4I4029/$1I2637/$1I43/MD ),
    .O(\$4I4029/$1I2637/Q0 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \$4I4029/$1I2637/$1I43/$1I32  (
    .I0(\$4I4029/$1I2637/$1N20 ),
    .I1(\$4I4029/$1I2637/Q0 ),
    .O(\$4I4029/$1I2637/$1I43/TQ )
  );
  X_AND2   \$4I4029/$1I2637/$1I43/$1I30/$1I9  (
    .I0(\$4I4029/$1I2637/$1N45 ),
    .I1(\$4I4029/$1I2637/$1N48 ),
    .O(\$4I4029/$1I2637/$1I43/$1I30/M1 )
  );
  X_OR2   \$4I4029/$1I2637/$1I43/$1I30/$1I8  (
    .I0(\$4I4029/$1I2637/$1I43/$1I30/M1 ),
    .I1(\$4I4029/$1I2637/$1I43/$1I30/M0 ),
    .O(\$4I4029/$1I2637/$1I43/MD )
  );
  X_AND2   \$4I4029/$1I2637/$1I43/$1I30/$1I7  (
    .I0(\NlwInverterSignal_$4I4029/$1I2637/$1I43/$1I30/$1I7/I0 ),
    .I1(\$4I4029/$1I2637/$1I43/TQ ),
    .O(\$4I4029/$1I2637/$1I43/$1I30/M0 )
  );
  X_ZERO   \$4I4029/$1I2637/$1I44/$1I2218  (
    .O(\$4I4029/$1I2637/$1I44/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2637/$1I44/L  (
    .I(\$4I4029/$1I2637/$1I44/$1N2216 ),
    .O(\$4I4029/$1I2637/$1N45 )
  );
  X_ZERO   \$4I4029/$1I2637/$1I47/$1I2218  (
    .O(\$4I4029/$1I2637/$1I47/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2637/$1I47/L  (
    .I(\$4I4029/$1I2637/$1I47/$1N2216 ),
    .O(\$4I4029/$1I2637/$1N48 )
  );
  X_ZERO   \$4I4029/$1I2637/$1I49/$1I2218  (
    .O(\$4I4029/$1I2637/$1I49/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2637/$1I49/L  (
    .I(\$4I4029/$1I2637/$1I49/$1N2216 ),
    .O(\$4I4029/$1I2637/$1N50 )
  );
  X_ZERO   \$4I4029/$1I2637/$1I52/$1I2218  (
    .O(\$4I4029/$1I2637/$1I52/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2637/$1I52/L  (
    .I(\$4I4029/$1I2637/$1I52/$1N2216 ),
    .O(\$4I4029/$1I2637/$1N51 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \$4I4029/$1I2637/$1I53/$1I35  (
    .CE(\$4I4029/$1N2734 ),
    .CLK(CLK),
    .I(\$4I4029/$1I2637/$1I53/MD ),
    .O(\$4I4029/$1I2637/Q1 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \$4I4029/$1I2637/$1I53/$1I32  (
    .I0(\$4I4029/$1I2637/Q0 ),
    .I1(\$4I4029/$1I2637/Q1 ),
    .O(\$4I4029/$1I2637/$1I53/TQ )
  );
  X_AND2   \$4I4029/$1I2637/$1I53/$1I30/$1I9  (
    .I0(\$4I4029/$1I2637/$1N50 ),
    .I1(\$4I4029/$1I2637/$1N51 ),
    .O(\$4I4029/$1I2637/$1I53/$1I30/M1 )
  );
  X_OR2   \$4I4029/$1I2637/$1I53/$1I30/$1I8  (
    .I0(\$4I4029/$1I2637/$1I53/$1I30/M1 ),
    .I1(\$4I4029/$1I2637/$1I53/$1I30/M0 ),
    .O(\$4I4029/$1I2637/$1I53/MD )
  );
  X_AND2   \$4I4029/$1I2637/$1I53/$1I30/$1I7  (
    .I0(\NlwInverterSignal_$4I4029/$1I2637/$1I53/$1I30/$1I7/I0 ),
    .I1(\$4I4029/$1I2637/$1I53/TQ ),
    .O(\$4I4029/$1I2637/$1I53/$1I30/M0 )
  );
  X_ZERO   \$4I4029/$1I2637/$1I54/$1I2218  (
    .O(\$4I4029/$1I2637/$1I54/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2637/$1I54/L  (
    .I(\$4I4029/$1I2637/$1I54/$1N2216 ),
    .O(\$4I4029/$1I2637/$1N55 )
  );
  X_ZERO   \$4I4029/$1I2637/$1I57/$1I2218  (
    .O(\$4I4029/$1I2637/$1I57/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2637/$1I57/L  (
    .I(\$4I4029/$1I2637/$1I57/$1N2216 ),
    .O(\$4I4029/$1I2637/$1N56 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \$4I4029/$1I2637/$1I58/$1I35  (
    .CE(\$4I4029/$1N2734 ),
    .CLK(CLK),
    .I(\$4I4029/$1I2637/$1I58/MD ),
    .O(\$4I4029/$1I2637/Q2 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \$4I4029/$1I2637/$1I58/$1I32  (
    .I0(\$4I4029/$1I2637/T2 ),
    .I1(\$4I4029/$1I2637/Q2 ),
    .O(\$4I4029/$1I2637/$1I58/TQ )
  );
  X_AND2   \$4I4029/$1I2637/$1I58/$1I30/$1I9  (
    .I0(\$4I4029/$1I2637/$1N55 ),
    .I1(\$4I4029/$1I2637/$1N56 ),
    .O(\$4I4029/$1I2637/$1I58/$1I30/M1 )
  );
  X_OR2   \$4I4029/$1I2637/$1I58/$1I30/$1I8  (
    .I0(\$4I4029/$1I2637/$1I58/$1I30/M1 ),
    .I1(\$4I4029/$1I2637/$1I58/$1I30/M0 ),
    .O(\$4I4029/$1I2637/$1I58/MD )
  );
  X_AND2   \$4I4029/$1I2637/$1I58/$1I30/$1I7  (
    .I0(\NlwInverterSignal_$4I4029/$1I2637/$1I58/$1I30/$1I7/I0 ),
    .I1(\$4I4029/$1I2637/$1I58/TQ ),
    .O(\$4I4029/$1I2637/$1I58/$1I30/M0 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \$4I4029/$1I2637/$1I59/$1I35  (
    .CE(\$4I4029/$1N2734 ),
    .CLK(CLK),
    .I(\$4I4029/$1I2637/$1I59/MD ),
    .O(\$4I4029/$1I2637/Q3 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \$4I4029/$1I2637/$1I59/$1I32  (
    .I0(\$4I4029/$1I2637/T3 ),
    .I1(\$4I4029/$1I2637/Q3 ),
    .O(\$4I4029/$1I2637/$1I59/TQ )
  );
  X_AND2   \$4I4029/$1I2637/$1I59/$1I30/$1I9  (
    .I0(\$4I4029/$1I2637/$1N62 ),
    .I1(\$4I4029/$1I2637/$1N61 ),
    .O(\$4I4029/$1I2637/$1I59/$1I30/M1 )
  );
  X_OR2   \$4I4029/$1I2637/$1I59/$1I30/$1I8  (
    .I0(\$4I4029/$1I2637/$1I59/$1I30/M1 ),
    .I1(\$4I4029/$1I2637/$1I59/$1I30/M0 ),
    .O(\$4I4029/$1I2637/$1I59/MD )
  );
  X_AND2   \$4I4029/$1I2637/$1I59/$1I30/$1I7  (
    .I0(\NlwInverterSignal_$4I4029/$1I2637/$1I59/$1I30/$1I7/I0 ),
    .I1(\$4I4029/$1I2637/$1I59/TQ ),
    .O(\$4I4029/$1I2637/$1I59/$1I30/M0 )
  );
  X_ZERO   \$4I4029/$1I2637/$1I60/$1I2218  (
    .O(\$4I4029/$1I2637/$1I60/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2637/$1I60/L  (
    .I(\$4I4029/$1I2637/$1I60/$1N2216 ),
    .O(\$4I4029/$1I2637/$1N61 )
  );
  X_ZERO   \$4I4029/$1I2637/$1I63/$1I2218  (
    .O(\$4I4029/$1I2637/$1I63/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2637/$1I63/L  (
    .I(\$4I4029/$1I2637/$1I63/$1N2216 ),
    .O(\$4I4029/$1I2637/$1N62 )
  );
  X_ZERO   \$4I4029/$1I2637/$1I64/$1I2218  (
    .O(\$4I4029/$1I2637/$1I64/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2637/$1I64/L  (
    .I(\$4I4029/$1I2637/$1I64/$1N2216 ),
    .O(\$4I4029/$1I2637/$1N65 )
  );
  X_ZERO   \$4I4029/$1I2637/$1I67/$1I2218  (
    .O(\$4I4029/$1I2637/$1I67/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2637/$1I67/L  (
    .I(\$4I4029/$1I2637/$1I67/$1N2216 ),
    .O(\$4I4029/$1I2637/$1N66 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \$4I4029/$1I2637/$1I68/$1I35  (
    .CE(\$4I4029/$1N2734 ),
    .CLK(CLK),
    .I(\$4I4029/$1I2637/$1I68/MD ),
    .O(\$4I4029/$1I2637/Q4 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \$4I4029/$1I2637/$1I68/$1I32  (
    .I0(\$4I4029/$1I2637/T4 ),
    .I1(\$4I4029/$1I2637/Q4 ),
    .O(\$4I4029/$1I2637/$1I68/TQ )
  );
  X_AND2   \$4I4029/$1I2637/$1I68/$1I30/$1I9  (
    .I0(\$4I4029/$1I2637/$1N65 ),
    .I1(\$4I4029/$1I2637/$1N66 ),
    .O(\$4I4029/$1I2637/$1I68/$1I30/M1 )
  );
  X_OR2   \$4I4029/$1I2637/$1I68/$1I30/$1I8  (
    .I0(\$4I4029/$1I2637/$1I68/$1I30/M1 ),
    .I1(\$4I4029/$1I2637/$1I68/$1I30/M0 ),
    .O(\$4I4029/$1I2637/$1I68/MD )
  );
  X_AND2   \$4I4029/$1I2637/$1I68/$1I30/$1I7  (
    .I0(\NlwInverterSignal_$4I4029/$1I2637/$1I68/$1I30/$1I7/I0 ),
    .I1(\$4I4029/$1I2637/$1I68/TQ ),
    .O(\$4I4029/$1I2637/$1I68/$1I30/M0 )
  );
  X_ZERO   \$4I4029/$1I2637/$1I69/$1I2218  (
    .O(\$4I4029/$1I2637/$1I69/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2637/$1I69/L  (
    .I(\$4I4029/$1I2637/$1I69/$1N2216 ),
    .O(\$4I4029/$1I2637/$1N70 )
  );
  X_ZERO   \$4I4029/$1I2637/$1I72/$1I2218  (
    .O(\$4I4029/$1I2637/$1I72/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2637/$1I72/L  (
    .I(\$4I4029/$1I2637/$1I72/$1N2216 ),
    .O(\$4I4029/$1I2637/$1N71 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \$4I4029/$1I2637/$1I73/$1I35  (
    .CE(\$4I4029/$1N2734 ),
    .CLK(CLK),
    .I(\$4I4029/$1I2637/$1I73/MD ),
    .O(\$4I4029/$1I2637/Q5 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \$4I4029/$1I2637/$1I73/$1I32  (
    .I0(\$4I4029/$1I2637/T5 ),
    .I1(\$4I4029/$1I2637/Q5 ),
    .O(\$4I4029/$1I2637/$1I73/TQ )
  );
  X_AND2   \$4I4029/$1I2637/$1I73/$1I30/$1I9  (
    .I0(\$4I4029/$1I2637/$1N70 ),
    .I1(\$4I4029/$1I2637/$1N71 ),
    .O(\$4I4029/$1I2637/$1I73/$1I30/M1 )
  );
  X_OR2   \$4I4029/$1I2637/$1I73/$1I30/$1I8  (
    .I0(\$4I4029/$1I2637/$1I73/$1I30/M1 ),
    .I1(\$4I4029/$1I2637/$1I73/$1I30/M0 ),
    .O(\$4I4029/$1I2637/$1I73/MD )
  );
  X_AND2   \$4I4029/$1I2637/$1I73/$1I30/$1I7  (
    .I0(\NlwInverterSignal_$4I4029/$1I2637/$1I73/$1I30/$1I7/I0 ),
    .I1(\$4I4029/$1I2637/$1I73/TQ ),
    .O(\$4I4029/$1I2637/$1I73/$1I30/M0 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \$4I4029/$1I2637/$1I79/$1I35  (
    .CE(\$4I4029/$1N2734 ),
    .CLK(CLK),
    .I(\$4I4029/$1I2637/$1I79/MD ),
    .O(\$4I4029/$1I2637/Q6 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \$4I4029/$1I2637/$1I79/$1I32  (
    .I0(\$4I4029/$1I2637/T6 ),
    .I1(\$4I4029/$1I2637/Q6 ),
    .O(\$4I4029/$1I2637/$1I79/TQ )
  );
  X_AND2   \$4I4029/$1I2637/$1I79/$1I30/$1I9  (
    .I0(\$4I4029/$1I2637/$1N82 ),
    .I1(\$4I4029/$1I2637/$1N81 ),
    .O(\$4I4029/$1I2637/$1I79/$1I30/M1 )
  );
  X_OR2   \$4I4029/$1I2637/$1I79/$1I30/$1I8  (
    .I0(\$4I4029/$1I2637/$1I79/$1I30/M1 ),
    .I1(\$4I4029/$1I2637/$1I79/$1I30/M0 ),
    .O(\$4I4029/$1I2637/$1I79/MD )
  );
  X_AND2   \$4I4029/$1I2637/$1I79/$1I30/$1I7  (
    .I0(\NlwInverterSignal_$4I4029/$1I2637/$1I79/$1I30/$1I7/I0 ),
    .I1(\$4I4029/$1I2637/$1I79/TQ ),
    .O(\$4I4029/$1I2637/$1I79/$1I30/M0 )
  );
  X_ZERO   \$4I4029/$1I2637/$1I80/$1I2218  (
    .O(\$4I4029/$1I2637/$1I80/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2637/$1I80/L  (
    .I(\$4I4029/$1I2637/$1I80/$1N2216 ),
    .O(\$4I4029/$1I2637/$1N81 )
  );
  X_ZERO   \$4I4029/$1I2637/$1I83/$1I2218  (
    .O(\$4I4029/$1I2637/$1I83/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2637/$1I83/L  (
    .I(\$4I4029/$1I2637/$1I83/$1N2216 ),
    .O(\$4I4029/$1I2637/$1N82 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \$4I4029/$1I2637/$1I84/$1I35  (
    .CE(\$4I4029/$1N2734 ),
    .CLK(CLK),
    .I(\$4I4029/$1I2637/$1I84/MD ),
    .O(\$4I4029/$1I2637/Q7 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \$4I4029/$1I2637/$1I84/$1I32  (
    .I0(\$4I4029/$1I2637/T7 ),
    .I1(\$4I4029/$1I2637/Q7 ),
    .O(\$4I4029/$1I2637/$1I84/TQ )
  );
  X_AND2   \$4I4029/$1I2637/$1I84/$1I30/$1I9  (
    .I0(\$4I4029/$1I2637/$1N87 ),
    .I1(\$4I4029/$1I2637/$1N86 ),
    .O(\$4I4029/$1I2637/$1I84/$1I30/M1 )
  );
  X_OR2   \$4I4029/$1I2637/$1I84/$1I30/$1I8  (
    .I0(\$4I4029/$1I2637/$1I84/$1I30/M1 ),
    .I1(\$4I4029/$1I2637/$1I84/$1I30/M0 ),
    .O(\$4I4029/$1I2637/$1I84/MD )
  );
  X_AND2   \$4I4029/$1I2637/$1I84/$1I30/$1I7  (
    .I0(\NlwInverterSignal_$4I4029/$1I2637/$1I84/$1I30/$1I7/I0 ),
    .I1(\$4I4029/$1I2637/$1I84/TQ ),
    .O(\$4I4029/$1I2637/$1I84/$1I30/M0 )
  );
  X_ZERO   \$4I4029/$1I2637/$1I85/$1I2218  (
    .O(\$4I4029/$1I2637/$1I85/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2637/$1I85/L  (
    .I(\$4I4029/$1I2637/$1I85/$1N2216 ),
    .O(\$4I4029/$1I2637/$1N86 )
  );
  X_ZERO   \$4I4029/$1I2637/$1I88/$1I2218  (
    .O(\$4I4029/$1I2637/$1I88/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2637/$1I88/L  (
    .I(\$4I4029/$1I2637/$1I88/$1N2216 ),
    .O(\$4I4029/$1I2637/$1N87 )
  );
  X_AND2   \$4I4029/$1I2645/$1I31  (
    .I0(\$4I4029/$1N2751 ),
    .I1(\$4I4029/$1I2645/TC ),
    .O(\$4I4029/$1N2753 )
  );
  X_AND4   \$4I4029/$1I2645/$1I28  (
    .I0(\$4I4029/$1I2645/Q6 ),
    .I1(\$4I4029/$1I2645/Q5 ),
    .I2(\$4I4029/$1I2645/Q4 ),
    .I3(\$4I4029/$1I2645/T4 ),
    .O(\$4I4029/$1I2645/T7 )
  );
  X_AND3   \$4I4029/$1I2645/$1I26  (
    .I0(\$4I4029/$1I2645/Q2 ),
    .I1(\$4I4029/$1I2645/Q1 ),
    .I2(\$4I4029/$1I2645/Q0 ),
    .O(\$4I4029/$1I2645/T3 )
  );
  X_AND2   \$4I4029/$1I2645/$1I24  (
    .I0(\$4I4029/$1I2645/Q1 ),
    .I1(\$4I4029/$1I2645/Q0 ),
    .O(\$4I4029/$1I2645/T2 )
  );
  X_AND2   \$4I4029/$1I2645/$1I2  (
    .I0(\$4I4029/$1I2645/Q4 ),
    .I1(\$4I4029/$1I2645/T4 ),
    .O(\$4I4029/$1I2645/T5 )
  );
  X_ONE   \$4I4029/$1I2645/$1I16  (
    .O(\$4I4029/$1I2645/$1N20 )
  );
  X_AND4   \$4I4029/$1I2645/$1I15  (
    .I0(\$4I4029/$1I2645/Q3 ),
    .I1(\$4I4029/$1I2645/Q2 ),
    .I2(\$4I4029/$1I2645/Q1 ),
    .I3(\$4I4029/$1I2645/Q0 ),
    .O(\$4I4029/$1I2645/T4 )
  );
  X_AND3   \$4I4029/$1I2645/$1I11  (
    .I0(\$4I4029/$1I2645/Q5 ),
    .I1(\$4I4029/$1I2645/Q4 ),
    .I2(\$4I4029/$1I2645/T4 ),
    .O(\$4I4029/$1I2645/T6 )
  );
  X_AND5   \$4I4029/$1I2645/$1I1  (
    .I0(\$4I4029/$1I2645/Q7 ),
    .I1(\$4I4029/$1I2645/Q6 ),
    .I2(\$4I4029/$1I2645/Q5 ),
    .I3(\$4I4029/$1I2645/Q4 ),
    .I4(\$4I4029/$1I2645/T4 ),
    .O(\$4I4029/$1I2645/TC )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \$4I4029/$1I2645/$1I43/$1I35  (
    .CE(\$4I4029/$1N2751 ),
    .CLK(CLK),
    .I(\$4I4029/$1I2645/$1I43/MD ),
    .O(\$4I4029/$1I2645/Q0 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \$4I4029/$1I2645/$1I43/$1I32  (
    .I0(\$4I4029/$1I2645/$1N20 ),
    .I1(\$4I4029/$1I2645/Q0 ),
    .O(\$4I4029/$1I2645/$1I43/TQ )
  );
  X_AND2   \$4I4029/$1I2645/$1I43/$1I30/$1I9  (
    .I0(\$4I4029/$1I2645/$1N45 ),
    .I1(\$4I4029/$1I2645/$1N48 ),
    .O(\$4I4029/$1I2645/$1I43/$1I30/M1 )
  );
  X_OR2   \$4I4029/$1I2645/$1I43/$1I30/$1I8  (
    .I0(\$4I4029/$1I2645/$1I43/$1I30/M1 ),
    .I1(\$4I4029/$1I2645/$1I43/$1I30/M0 ),
    .O(\$4I4029/$1I2645/$1I43/MD )
  );
  X_AND2   \$4I4029/$1I2645/$1I43/$1I30/$1I7  (
    .I0(\NlwInverterSignal_$4I4029/$1I2645/$1I43/$1I30/$1I7/I0 ),
    .I1(\$4I4029/$1I2645/$1I43/TQ ),
    .O(\$4I4029/$1I2645/$1I43/$1I30/M0 )
  );
  X_ZERO   \$4I4029/$1I2645/$1I44/$1I2218  (
    .O(\$4I4029/$1I2645/$1I44/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2645/$1I44/L  (
    .I(\$4I4029/$1I2645/$1I44/$1N2216 ),
    .O(\$4I4029/$1I2645/$1N45 )
  );
  X_ZERO   \$4I4029/$1I2645/$1I47/$1I2218  (
    .O(\$4I4029/$1I2645/$1I47/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2645/$1I47/L  (
    .I(\$4I4029/$1I2645/$1I47/$1N2216 ),
    .O(\$4I4029/$1I2645/$1N48 )
  );
  X_ZERO   \$4I4029/$1I2645/$1I49/$1I2218  (
    .O(\$4I4029/$1I2645/$1I49/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2645/$1I49/L  (
    .I(\$4I4029/$1I2645/$1I49/$1N2216 ),
    .O(\$4I4029/$1I2645/$1N50 )
  );
  X_ZERO   \$4I4029/$1I2645/$1I52/$1I2218  (
    .O(\$4I4029/$1I2645/$1I52/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2645/$1I52/L  (
    .I(\$4I4029/$1I2645/$1I52/$1N2216 ),
    .O(\$4I4029/$1I2645/$1N51 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \$4I4029/$1I2645/$1I53/$1I35  (
    .CE(\$4I4029/$1N2751 ),
    .CLK(CLK),
    .I(\$4I4029/$1I2645/$1I53/MD ),
    .O(\$4I4029/$1I2645/Q1 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \$4I4029/$1I2645/$1I53/$1I32  (
    .I0(\$4I4029/$1I2645/Q0 ),
    .I1(\$4I4029/$1I2645/Q1 ),
    .O(\$4I4029/$1I2645/$1I53/TQ )
  );
  X_AND2   \$4I4029/$1I2645/$1I53/$1I30/$1I9  (
    .I0(\$4I4029/$1I2645/$1N50 ),
    .I1(\$4I4029/$1I2645/$1N51 ),
    .O(\$4I4029/$1I2645/$1I53/$1I30/M1 )
  );
  X_OR2   \$4I4029/$1I2645/$1I53/$1I30/$1I8  (
    .I0(\$4I4029/$1I2645/$1I53/$1I30/M1 ),
    .I1(\$4I4029/$1I2645/$1I53/$1I30/M0 ),
    .O(\$4I4029/$1I2645/$1I53/MD )
  );
  X_AND2   \$4I4029/$1I2645/$1I53/$1I30/$1I7  (
    .I0(\NlwInverterSignal_$4I4029/$1I2645/$1I53/$1I30/$1I7/I0 ),
    .I1(\$4I4029/$1I2645/$1I53/TQ ),
    .O(\$4I4029/$1I2645/$1I53/$1I30/M0 )
  );
  X_ZERO   \$4I4029/$1I2645/$1I54/$1I2218  (
    .O(\$4I4029/$1I2645/$1I54/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2645/$1I54/L  (
    .I(\$4I4029/$1I2645/$1I54/$1N2216 ),
    .O(\$4I4029/$1I2645/$1N55 )
  );
  X_ZERO   \$4I4029/$1I2645/$1I57/$1I2218  (
    .O(\$4I4029/$1I2645/$1I57/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2645/$1I57/L  (
    .I(\$4I4029/$1I2645/$1I57/$1N2216 ),
    .O(\$4I4029/$1I2645/$1N56 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \$4I4029/$1I2645/$1I58/$1I35  (
    .CE(\$4I4029/$1N2751 ),
    .CLK(CLK),
    .I(\$4I4029/$1I2645/$1I58/MD ),
    .O(\$4I4029/$1I2645/Q2 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \$4I4029/$1I2645/$1I58/$1I32  (
    .I0(\$4I4029/$1I2645/T2 ),
    .I1(\$4I4029/$1I2645/Q2 ),
    .O(\$4I4029/$1I2645/$1I58/TQ )
  );
  X_AND2   \$4I4029/$1I2645/$1I58/$1I30/$1I9  (
    .I0(\$4I4029/$1I2645/$1N55 ),
    .I1(\$4I4029/$1I2645/$1N56 ),
    .O(\$4I4029/$1I2645/$1I58/$1I30/M1 )
  );
  X_OR2   \$4I4029/$1I2645/$1I58/$1I30/$1I8  (
    .I0(\$4I4029/$1I2645/$1I58/$1I30/M1 ),
    .I1(\$4I4029/$1I2645/$1I58/$1I30/M0 ),
    .O(\$4I4029/$1I2645/$1I58/MD )
  );
  X_AND2   \$4I4029/$1I2645/$1I58/$1I30/$1I7  (
    .I0(\NlwInverterSignal_$4I4029/$1I2645/$1I58/$1I30/$1I7/I0 ),
    .I1(\$4I4029/$1I2645/$1I58/TQ ),
    .O(\$4I4029/$1I2645/$1I58/$1I30/M0 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \$4I4029/$1I2645/$1I59/$1I35  (
    .CE(\$4I4029/$1N2751 ),
    .CLK(CLK),
    .I(\$4I4029/$1I2645/$1I59/MD ),
    .O(\$4I4029/$1I2645/Q3 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \$4I4029/$1I2645/$1I59/$1I32  (
    .I0(\$4I4029/$1I2645/T3 ),
    .I1(\$4I4029/$1I2645/Q3 ),
    .O(\$4I4029/$1I2645/$1I59/TQ )
  );
  X_AND2   \$4I4029/$1I2645/$1I59/$1I30/$1I9  (
    .I0(\$4I4029/$1I2645/$1N62 ),
    .I1(\$4I4029/$1I2645/$1N61 ),
    .O(\$4I4029/$1I2645/$1I59/$1I30/M1 )
  );
  X_OR2   \$4I4029/$1I2645/$1I59/$1I30/$1I8  (
    .I0(\$4I4029/$1I2645/$1I59/$1I30/M1 ),
    .I1(\$4I4029/$1I2645/$1I59/$1I30/M0 ),
    .O(\$4I4029/$1I2645/$1I59/MD )
  );
  X_AND2   \$4I4029/$1I2645/$1I59/$1I30/$1I7  (
    .I0(\NlwInverterSignal_$4I4029/$1I2645/$1I59/$1I30/$1I7/I0 ),
    .I1(\$4I4029/$1I2645/$1I59/TQ ),
    .O(\$4I4029/$1I2645/$1I59/$1I30/M0 )
  );
  X_ZERO   \$4I4029/$1I2645/$1I60/$1I2218  (
    .O(\$4I4029/$1I2645/$1I60/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2645/$1I60/L  (
    .I(\$4I4029/$1I2645/$1I60/$1N2216 ),
    .O(\$4I4029/$1I2645/$1N61 )
  );
  X_ZERO   \$4I4029/$1I2645/$1I63/$1I2218  (
    .O(\$4I4029/$1I2645/$1I63/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2645/$1I63/L  (
    .I(\$4I4029/$1I2645/$1I63/$1N2216 ),
    .O(\$4I4029/$1I2645/$1N62 )
  );
  X_ZERO   \$4I4029/$1I2645/$1I64/$1I2218  (
    .O(\$4I4029/$1I2645/$1I64/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2645/$1I64/L  (
    .I(\$4I4029/$1I2645/$1I64/$1N2216 ),
    .O(\$4I4029/$1I2645/$1N65 )
  );
  X_ZERO   \$4I4029/$1I2645/$1I67/$1I2218  (
    .O(\$4I4029/$1I2645/$1I67/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2645/$1I67/L  (
    .I(\$4I4029/$1I2645/$1I67/$1N2216 ),
    .O(\$4I4029/$1I2645/$1N66 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \$4I4029/$1I2645/$1I68/$1I35  (
    .CE(\$4I4029/$1N2751 ),
    .CLK(CLK),
    .I(\$4I4029/$1I2645/$1I68/MD ),
    .O(\$4I4029/$1I2645/Q4 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \$4I4029/$1I2645/$1I68/$1I32  (
    .I0(\$4I4029/$1I2645/T4 ),
    .I1(\$4I4029/$1I2645/Q4 ),
    .O(\$4I4029/$1I2645/$1I68/TQ )
  );
  X_AND2   \$4I4029/$1I2645/$1I68/$1I30/$1I9  (
    .I0(\$4I4029/$1I2645/$1N65 ),
    .I1(\$4I4029/$1I2645/$1N66 ),
    .O(\$4I4029/$1I2645/$1I68/$1I30/M1 )
  );
  X_OR2   \$4I4029/$1I2645/$1I68/$1I30/$1I8  (
    .I0(\$4I4029/$1I2645/$1I68/$1I30/M1 ),
    .I1(\$4I4029/$1I2645/$1I68/$1I30/M0 ),
    .O(\$4I4029/$1I2645/$1I68/MD )
  );
  X_AND2   \$4I4029/$1I2645/$1I68/$1I30/$1I7  (
    .I0(\NlwInverterSignal_$4I4029/$1I2645/$1I68/$1I30/$1I7/I0 ),
    .I1(\$4I4029/$1I2645/$1I68/TQ ),
    .O(\$4I4029/$1I2645/$1I68/$1I30/M0 )
  );
  X_ZERO   \$4I4029/$1I2645/$1I69/$1I2218  (
    .O(\$4I4029/$1I2645/$1I69/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2645/$1I69/L  (
    .I(\$4I4029/$1I2645/$1I69/$1N2216 ),
    .O(\$4I4029/$1I2645/$1N70 )
  );
  X_ZERO   \$4I4029/$1I2645/$1I72/$1I2218  (
    .O(\$4I4029/$1I2645/$1I72/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2645/$1I72/L  (
    .I(\$4I4029/$1I2645/$1I72/$1N2216 ),
    .O(\$4I4029/$1I2645/$1N71 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \$4I4029/$1I2645/$1I73/$1I35  (
    .CE(\$4I4029/$1N2751 ),
    .CLK(CLK),
    .I(\$4I4029/$1I2645/$1I73/MD ),
    .O(\$4I4029/$1I2645/Q5 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \$4I4029/$1I2645/$1I73/$1I32  (
    .I0(\$4I4029/$1I2645/T5 ),
    .I1(\$4I4029/$1I2645/Q5 ),
    .O(\$4I4029/$1I2645/$1I73/TQ )
  );
  X_AND2   \$4I4029/$1I2645/$1I73/$1I30/$1I9  (
    .I0(\$4I4029/$1I2645/$1N70 ),
    .I1(\$4I4029/$1I2645/$1N71 ),
    .O(\$4I4029/$1I2645/$1I73/$1I30/M1 )
  );
  X_OR2   \$4I4029/$1I2645/$1I73/$1I30/$1I8  (
    .I0(\$4I4029/$1I2645/$1I73/$1I30/M1 ),
    .I1(\$4I4029/$1I2645/$1I73/$1I30/M0 ),
    .O(\$4I4029/$1I2645/$1I73/MD )
  );
  X_AND2   \$4I4029/$1I2645/$1I73/$1I30/$1I7  (
    .I0(\NlwInverterSignal_$4I4029/$1I2645/$1I73/$1I30/$1I7/I0 ),
    .I1(\$4I4029/$1I2645/$1I73/TQ ),
    .O(\$4I4029/$1I2645/$1I73/$1I30/M0 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \$4I4029/$1I2645/$1I79/$1I35  (
    .CE(\$4I4029/$1N2751 ),
    .CLK(CLK),
    .I(\$4I4029/$1I2645/$1I79/MD ),
    .O(\$4I4029/$1I2645/Q6 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \$4I4029/$1I2645/$1I79/$1I32  (
    .I0(\$4I4029/$1I2645/T6 ),
    .I1(\$4I4029/$1I2645/Q6 ),
    .O(\$4I4029/$1I2645/$1I79/TQ )
  );
  X_AND2   \$4I4029/$1I2645/$1I79/$1I30/$1I9  (
    .I0(\$4I4029/$1I2645/$1N82 ),
    .I1(\$4I4029/$1I2645/$1N81 ),
    .O(\$4I4029/$1I2645/$1I79/$1I30/M1 )
  );
  X_OR2   \$4I4029/$1I2645/$1I79/$1I30/$1I8  (
    .I0(\$4I4029/$1I2645/$1I79/$1I30/M1 ),
    .I1(\$4I4029/$1I2645/$1I79/$1I30/M0 ),
    .O(\$4I4029/$1I2645/$1I79/MD )
  );
  X_AND2   \$4I4029/$1I2645/$1I79/$1I30/$1I7  (
    .I0(\NlwInverterSignal_$4I4029/$1I2645/$1I79/$1I30/$1I7/I0 ),
    .I1(\$4I4029/$1I2645/$1I79/TQ ),
    .O(\$4I4029/$1I2645/$1I79/$1I30/M0 )
  );
  X_ZERO   \$4I4029/$1I2645/$1I80/$1I2218  (
    .O(\$4I4029/$1I2645/$1I80/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2645/$1I80/L  (
    .I(\$4I4029/$1I2645/$1I80/$1N2216 ),
    .O(\$4I4029/$1I2645/$1N81 )
  );
  X_ZERO   \$4I4029/$1I2645/$1I83/$1I2218  (
    .O(\$4I4029/$1I2645/$1I83/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2645/$1I83/L  (
    .I(\$4I4029/$1I2645/$1I83/$1N2216 ),
    .O(\$4I4029/$1I2645/$1N82 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \$4I4029/$1I2645/$1I84/$1I35  (
    .CE(\$4I4029/$1N2751 ),
    .CLK(CLK),
    .I(\$4I4029/$1I2645/$1I84/MD ),
    .O(\$4I4029/$1I2645/Q7 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \$4I4029/$1I2645/$1I84/$1I32  (
    .I0(\$4I4029/$1I2645/T7 ),
    .I1(\$4I4029/$1I2645/Q7 ),
    .O(\$4I4029/$1I2645/$1I84/TQ )
  );
  X_AND2   \$4I4029/$1I2645/$1I84/$1I30/$1I9  (
    .I0(\$4I4029/$1I2645/$1N87 ),
    .I1(\$4I4029/$1I2645/$1N86 ),
    .O(\$4I4029/$1I2645/$1I84/$1I30/M1 )
  );
  X_OR2   \$4I4029/$1I2645/$1I84/$1I30/$1I8  (
    .I0(\$4I4029/$1I2645/$1I84/$1I30/M1 ),
    .I1(\$4I4029/$1I2645/$1I84/$1I30/M0 ),
    .O(\$4I4029/$1I2645/$1I84/MD )
  );
  X_AND2   \$4I4029/$1I2645/$1I84/$1I30/$1I7  (
    .I0(\NlwInverterSignal_$4I4029/$1I2645/$1I84/$1I30/$1I7/I0 ),
    .I1(\$4I4029/$1I2645/$1I84/TQ ),
    .O(\$4I4029/$1I2645/$1I84/$1I30/M0 )
  );
  X_ZERO   \$4I4029/$1I2645/$1I85/$1I2218  (
    .O(\$4I4029/$1I2645/$1I85/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2645/$1I85/L  (
    .I(\$4I4029/$1I2645/$1I85/$1N2216 ),
    .O(\$4I4029/$1I2645/$1N86 )
  );
  X_ZERO   \$4I4029/$1I2645/$1I88/$1I2218  (
    .O(\$4I4029/$1I2645/$1I88/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2645/$1I88/L  (
    .I(\$4I4029/$1I2645/$1I88/$1N2216 ),
    .O(\$4I4029/$1I2645/$1N87 )
  );
  X_AND2   \$4I4029/$1I2653/$1I31  (
    .I0(\$4I4029/$1N2755 ),
    .I1(\$4I4029/$1I2653/TC ),
    .O(\$4I4029/$1N2757 )
  );
  X_AND4   \$4I4029/$1I2653/$1I28  (
    .I0(\$4I4029/$1I2653/Q6 ),
    .I1(\$4I4029/$1I2653/Q5 ),
    .I2(\$4I4029/$1I2653/Q4 ),
    .I3(\$4I4029/$1I2653/T4 ),
    .O(\$4I4029/$1I2653/T7 )
  );
  X_AND3   \$4I4029/$1I2653/$1I26  (
    .I0(\$4I4029/$1I2653/Q2 ),
    .I1(\$4I4029/$1I2653/Q1 ),
    .I2(\$4I4029/$1I2653/Q0 ),
    .O(\$4I4029/$1I2653/T3 )
  );
  X_AND2   \$4I4029/$1I2653/$1I24  (
    .I0(\$4I4029/$1I2653/Q1 ),
    .I1(\$4I4029/$1I2653/Q0 ),
    .O(\$4I4029/$1I2653/T2 )
  );
  X_AND2   \$4I4029/$1I2653/$1I2  (
    .I0(\$4I4029/$1I2653/Q4 ),
    .I1(\$4I4029/$1I2653/T4 ),
    .O(\$4I4029/$1I2653/T5 )
  );
  X_ONE   \$4I4029/$1I2653/$1I16  (
    .O(\$4I4029/$1I2653/$1N20 )
  );
  X_AND4   \$4I4029/$1I2653/$1I15  (
    .I0(\$4I4029/$1I2653/Q3 ),
    .I1(\$4I4029/$1I2653/Q2 ),
    .I2(\$4I4029/$1I2653/Q1 ),
    .I3(\$4I4029/$1I2653/Q0 ),
    .O(\$4I4029/$1I2653/T4 )
  );
  X_AND3   \$4I4029/$1I2653/$1I11  (
    .I0(\$4I4029/$1I2653/Q5 ),
    .I1(\$4I4029/$1I2653/Q4 ),
    .I2(\$4I4029/$1I2653/T4 ),
    .O(\$4I4029/$1I2653/T6 )
  );
  X_AND5   \$4I4029/$1I2653/$1I1  (
    .I0(\$4I4029/$1I2653/Q7 ),
    .I1(\$4I4029/$1I2653/Q6 ),
    .I2(\$4I4029/$1I2653/Q5 ),
    .I3(\$4I4029/$1I2653/Q4 ),
    .I4(\$4I4029/$1I2653/T4 ),
    .O(\$4I4029/$1I2653/TC )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \$4I4029/$1I2653/$1I43/$1I35  (
    .CE(\$4I4029/$1N2755 ),
    .CLK(CLK),
    .I(\$4I4029/$1I2653/$1I43/MD ),
    .O(\$4I4029/$1I2653/Q0 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \$4I4029/$1I2653/$1I43/$1I32  (
    .I0(\$4I4029/$1I2653/$1N20 ),
    .I1(\$4I4029/$1I2653/Q0 ),
    .O(\$4I4029/$1I2653/$1I43/TQ )
  );
  X_AND2   \$4I4029/$1I2653/$1I43/$1I30/$1I9  (
    .I0(\$4I4029/$1I2653/$1N45 ),
    .I1(\$4I4029/$1I2653/$1N48 ),
    .O(\$4I4029/$1I2653/$1I43/$1I30/M1 )
  );
  X_OR2   \$4I4029/$1I2653/$1I43/$1I30/$1I8  (
    .I0(\$4I4029/$1I2653/$1I43/$1I30/M1 ),
    .I1(\$4I4029/$1I2653/$1I43/$1I30/M0 ),
    .O(\$4I4029/$1I2653/$1I43/MD )
  );
  X_AND2   \$4I4029/$1I2653/$1I43/$1I30/$1I7  (
    .I0(\NlwInverterSignal_$4I4029/$1I2653/$1I43/$1I30/$1I7/I0 ),
    .I1(\$4I4029/$1I2653/$1I43/TQ ),
    .O(\$4I4029/$1I2653/$1I43/$1I30/M0 )
  );
  X_ZERO   \$4I4029/$1I2653/$1I44/$1I2218  (
    .O(\$4I4029/$1I2653/$1I44/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2653/$1I44/L  (
    .I(\$4I4029/$1I2653/$1I44/$1N2216 ),
    .O(\$4I4029/$1I2653/$1N45 )
  );
  X_ZERO   \$4I4029/$1I2653/$1I47/$1I2218  (
    .O(\$4I4029/$1I2653/$1I47/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2653/$1I47/L  (
    .I(\$4I4029/$1I2653/$1I47/$1N2216 ),
    .O(\$4I4029/$1I2653/$1N48 )
  );
  X_ZERO   \$4I4029/$1I2653/$1I49/$1I2218  (
    .O(\$4I4029/$1I2653/$1I49/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2653/$1I49/L  (
    .I(\$4I4029/$1I2653/$1I49/$1N2216 ),
    .O(\$4I4029/$1I2653/$1N50 )
  );
  X_ZERO   \$4I4029/$1I2653/$1I52/$1I2218  (
    .O(\$4I4029/$1I2653/$1I52/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2653/$1I52/L  (
    .I(\$4I4029/$1I2653/$1I52/$1N2216 ),
    .O(\$4I4029/$1I2653/$1N51 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \$4I4029/$1I2653/$1I53/$1I35  (
    .CE(\$4I4029/$1N2755 ),
    .CLK(CLK),
    .I(\$4I4029/$1I2653/$1I53/MD ),
    .O(\$4I4029/$1I2653/Q1 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \$4I4029/$1I2653/$1I53/$1I32  (
    .I0(\$4I4029/$1I2653/Q0 ),
    .I1(\$4I4029/$1I2653/Q1 ),
    .O(\$4I4029/$1I2653/$1I53/TQ )
  );
  X_AND2   \$4I4029/$1I2653/$1I53/$1I30/$1I9  (
    .I0(\$4I4029/$1I2653/$1N50 ),
    .I1(\$4I4029/$1I2653/$1N51 ),
    .O(\$4I4029/$1I2653/$1I53/$1I30/M1 )
  );
  X_OR2   \$4I4029/$1I2653/$1I53/$1I30/$1I8  (
    .I0(\$4I4029/$1I2653/$1I53/$1I30/M1 ),
    .I1(\$4I4029/$1I2653/$1I53/$1I30/M0 ),
    .O(\$4I4029/$1I2653/$1I53/MD )
  );
  X_AND2   \$4I4029/$1I2653/$1I53/$1I30/$1I7  (
    .I0(\NlwInverterSignal_$4I4029/$1I2653/$1I53/$1I30/$1I7/I0 ),
    .I1(\$4I4029/$1I2653/$1I53/TQ ),
    .O(\$4I4029/$1I2653/$1I53/$1I30/M0 )
  );
  X_ZERO   \$4I4029/$1I2653/$1I54/$1I2218  (
    .O(\$4I4029/$1I2653/$1I54/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2653/$1I54/L  (
    .I(\$4I4029/$1I2653/$1I54/$1N2216 ),
    .O(\$4I4029/$1I2653/$1N55 )
  );
  X_ZERO   \$4I4029/$1I2653/$1I57/$1I2218  (
    .O(\$4I4029/$1I2653/$1I57/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2653/$1I57/L  (
    .I(\$4I4029/$1I2653/$1I57/$1N2216 ),
    .O(\$4I4029/$1I2653/$1N56 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \$4I4029/$1I2653/$1I58/$1I35  (
    .CE(\$4I4029/$1N2755 ),
    .CLK(CLK),
    .I(\$4I4029/$1I2653/$1I58/MD ),
    .O(\$4I4029/$1I2653/Q2 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \$4I4029/$1I2653/$1I58/$1I32  (
    .I0(\$4I4029/$1I2653/T2 ),
    .I1(\$4I4029/$1I2653/Q2 ),
    .O(\$4I4029/$1I2653/$1I58/TQ )
  );
  X_AND2   \$4I4029/$1I2653/$1I58/$1I30/$1I9  (
    .I0(\$4I4029/$1I2653/$1N55 ),
    .I1(\$4I4029/$1I2653/$1N56 ),
    .O(\$4I4029/$1I2653/$1I58/$1I30/M1 )
  );
  X_OR2   \$4I4029/$1I2653/$1I58/$1I30/$1I8  (
    .I0(\$4I4029/$1I2653/$1I58/$1I30/M1 ),
    .I1(\$4I4029/$1I2653/$1I58/$1I30/M0 ),
    .O(\$4I4029/$1I2653/$1I58/MD )
  );
  X_AND2   \$4I4029/$1I2653/$1I58/$1I30/$1I7  (
    .I0(\NlwInverterSignal_$4I4029/$1I2653/$1I58/$1I30/$1I7/I0 ),
    .I1(\$4I4029/$1I2653/$1I58/TQ ),
    .O(\$4I4029/$1I2653/$1I58/$1I30/M0 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \$4I4029/$1I2653/$1I59/$1I35  (
    .CE(\$4I4029/$1N2755 ),
    .CLK(CLK),
    .I(\$4I4029/$1I2653/$1I59/MD ),
    .O(\$4I4029/$1I2653/Q3 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \$4I4029/$1I2653/$1I59/$1I32  (
    .I0(\$4I4029/$1I2653/T3 ),
    .I1(\$4I4029/$1I2653/Q3 ),
    .O(\$4I4029/$1I2653/$1I59/TQ )
  );
  X_AND2   \$4I4029/$1I2653/$1I59/$1I30/$1I9  (
    .I0(\$4I4029/$1I2653/$1N62 ),
    .I1(\$4I4029/$1I2653/$1N61 ),
    .O(\$4I4029/$1I2653/$1I59/$1I30/M1 )
  );
  X_OR2   \$4I4029/$1I2653/$1I59/$1I30/$1I8  (
    .I0(\$4I4029/$1I2653/$1I59/$1I30/M1 ),
    .I1(\$4I4029/$1I2653/$1I59/$1I30/M0 ),
    .O(\$4I4029/$1I2653/$1I59/MD )
  );
  X_AND2   \$4I4029/$1I2653/$1I59/$1I30/$1I7  (
    .I0(\NlwInverterSignal_$4I4029/$1I2653/$1I59/$1I30/$1I7/I0 ),
    .I1(\$4I4029/$1I2653/$1I59/TQ ),
    .O(\$4I4029/$1I2653/$1I59/$1I30/M0 )
  );
  X_ZERO   \$4I4029/$1I2653/$1I60/$1I2218  (
    .O(\$4I4029/$1I2653/$1I60/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2653/$1I60/L  (
    .I(\$4I4029/$1I2653/$1I60/$1N2216 ),
    .O(\$4I4029/$1I2653/$1N61 )
  );
  X_ZERO   \$4I4029/$1I2653/$1I63/$1I2218  (
    .O(\$4I4029/$1I2653/$1I63/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2653/$1I63/L  (
    .I(\$4I4029/$1I2653/$1I63/$1N2216 ),
    .O(\$4I4029/$1I2653/$1N62 )
  );
  X_ZERO   \$4I4029/$1I2653/$1I64/$1I2218  (
    .O(\$4I4029/$1I2653/$1I64/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2653/$1I64/L  (
    .I(\$4I4029/$1I2653/$1I64/$1N2216 ),
    .O(\$4I4029/$1I2653/$1N65 )
  );
  X_ZERO   \$4I4029/$1I2653/$1I67/$1I2218  (
    .O(\$4I4029/$1I2653/$1I67/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2653/$1I67/L  (
    .I(\$4I4029/$1I2653/$1I67/$1N2216 ),
    .O(\$4I4029/$1I2653/$1N66 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \$4I4029/$1I2653/$1I68/$1I35  (
    .CE(\$4I4029/$1N2755 ),
    .CLK(CLK),
    .I(\$4I4029/$1I2653/$1I68/MD ),
    .O(\$4I4029/$1I2653/Q4 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \$4I4029/$1I2653/$1I68/$1I32  (
    .I0(\$4I4029/$1I2653/T4 ),
    .I1(\$4I4029/$1I2653/Q4 ),
    .O(\$4I4029/$1I2653/$1I68/TQ )
  );
  X_AND2   \$4I4029/$1I2653/$1I68/$1I30/$1I9  (
    .I0(\$4I4029/$1I2653/$1N65 ),
    .I1(\$4I4029/$1I2653/$1N66 ),
    .O(\$4I4029/$1I2653/$1I68/$1I30/M1 )
  );
  X_OR2   \$4I4029/$1I2653/$1I68/$1I30/$1I8  (
    .I0(\$4I4029/$1I2653/$1I68/$1I30/M1 ),
    .I1(\$4I4029/$1I2653/$1I68/$1I30/M0 ),
    .O(\$4I4029/$1I2653/$1I68/MD )
  );
  X_AND2   \$4I4029/$1I2653/$1I68/$1I30/$1I7  (
    .I0(\NlwInverterSignal_$4I4029/$1I2653/$1I68/$1I30/$1I7/I0 ),
    .I1(\$4I4029/$1I2653/$1I68/TQ ),
    .O(\$4I4029/$1I2653/$1I68/$1I30/M0 )
  );
  X_ZERO   \$4I4029/$1I2653/$1I69/$1I2218  (
    .O(\$4I4029/$1I2653/$1I69/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2653/$1I69/L  (
    .I(\$4I4029/$1I2653/$1I69/$1N2216 ),
    .O(\$4I4029/$1I2653/$1N70 )
  );
  X_ZERO   \$4I4029/$1I2653/$1I72/$1I2218  (
    .O(\$4I4029/$1I2653/$1I72/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2653/$1I72/L  (
    .I(\$4I4029/$1I2653/$1I72/$1N2216 ),
    .O(\$4I4029/$1I2653/$1N71 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \$4I4029/$1I2653/$1I73/$1I35  (
    .CE(\$4I4029/$1N2755 ),
    .CLK(CLK),
    .I(\$4I4029/$1I2653/$1I73/MD ),
    .O(\$4I4029/$1I2653/Q5 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \$4I4029/$1I2653/$1I73/$1I32  (
    .I0(\$4I4029/$1I2653/T5 ),
    .I1(\$4I4029/$1I2653/Q5 ),
    .O(\$4I4029/$1I2653/$1I73/TQ )
  );
  X_AND2   \$4I4029/$1I2653/$1I73/$1I30/$1I9  (
    .I0(\$4I4029/$1I2653/$1N70 ),
    .I1(\$4I4029/$1I2653/$1N71 ),
    .O(\$4I4029/$1I2653/$1I73/$1I30/M1 )
  );
  X_OR2   \$4I4029/$1I2653/$1I73/$1I30/$1I8  (
    .I0(\$4I4029/$1I2653/$1I73/$1I30/M1 ),
    .I1(\$4I4029/$1I2653/$1I73/$1I30/M0 ),
    .O(\$4I4029/$1I2653/$1I73/MD )
  );
  X_AND2   \$4I4029/$1I2653/$1I73/$1I30/$1I7  (
    .I0(\NlwInverterSignal_$4I4029/$1I2653/$1I73/$1I30/$1I7/I0 ),
    .I1(\$4I4029/$1I2653/$1I73/TQ ),
    .O(\$4I4029/$1I2653/$1I73/$1I30/M0 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \$4I4029/$1I2653/$1I79/$1I35  (
    .CE(\$4I4029/$1N2755 ),
    .CLK(CLK),
    .I(\$4I4029/$1I2653/$1I79/MD ),
    .O(\$4I4029/$1I2653/Q6 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \$4I4029/$1I2653/$1I79/$1I32  (
    .I0(\$4I4029/$1I2653/T6 ),
    .I1(\$4I4029/$1I2653/Q6 ),
    .O(\$4I4029/$1I2653/$1I79/TQ )
  );
  X_AND2   \$4I4029/$1I2653/$1I79/$1I30/$1I9  (
    .I0(\$4I4029/$1I2653/$1N82 ),
    .I1(\$4I4029/$1I2653/$1N81 ),
    .O(\$4I4029/$1I2653/$1I79/$1I30/M1 )
  );
  X_OR2   \$4I4029/$1I2653/$1I79/$1I30/$1I8  (
    .I0(\$4I4029/$1I2653/$1I79/$1I30/M1 ),
    .I1(\$4I4029/$1I2653/$1I79/$1I30/M0 ),
    .O(\$4I4029/$1I2653/$1I79/MD )
  );
  X_AND2   \$4I4029/$1I2653/$1I79/$1I30/$1I7  (
    .I0(\NlwInverterSignal_$4I4029/$1I2653/$1I79/$1I30/$1I7/I0 ),
    .I1(\$4I4029/$1I2653/$1I79/TQ ),
    .O(\$4I4029/$1I2653/$1I79/$1I30/M0 )
  );
  X_ZERO   \$4I4029/$1I2653/$1I80/$1I2218  (
    .O(\$4I4029/$1I2653/$1I80/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2653/$1I80/L  (
    .I(\$4I4029/$1I2653/$1I80/$1N2216 ),
    .O(\$4I4029/$1I2653/$1N81 )
  );
  X_ZERO   \$4I4029/$1I2653/$1I83/$1I2218  (
    .O(\$4I4029/$1I2653/$1I83/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2653/$1I83/L  (
    .I(\$4I4029/$1I2653/$1I83/$1N2216 ),
    .O(\$4I4029/$1I2653/$1N82 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \$4I4029/$1I2653/$1I84/$1I35  (
    .CE(\$4I4029/$1N2755 ),
    .CLK(CLK),
    .I(\$4I4029/$1I2653/$1I84/MD ),
    .O(\$4I4029/$1I2653/Q7 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \$4I4029/$1I2653/$1I84/$1I32  (
    .I0(\$4I4029/$1I2653/T7 ),
    .I1(\$4I4029/$1I2653/Q7 ),
    .O(\$4I4029/$1I2653/$1I84/TQ )
  );
  X_AND2   \$4I4029/$1I2653/$1I84/$1I30/$1I9  (
    .I0(\$4I4029/$1I2653/$1N87 ),
    .I1(\$4I4029/$1I2653/$1N86 ),
    .O(\$4I4029/$1I2653/$1I84/$1I30/M1 )
  );
  X_OR2   \$4I4029/$1I2653/$1I84/$1I30/$1I8  (
    .I0(\$4I4029/$1I2653/$1I84/$1I30/M1 ),
    .I1(\$4I4029/$1I2653/$1I84/$1I30/M0 ),
    .O(\$4I4029/$1I2653/$1I84/MD )
  );
  X_AND2   \$4I4029/$1I2653/$1I84/$1I30/$1I7  (
    .I0(\NlwInverterSignal_$4I4029/$1I2653/$1I84/$1I30/$1I7/I0 ),
    .I1(\$4I4029/$1I2653/$1I84/TQ ),
    .O(\$4I4029/$1I2653/$1I84/$1I30/M0 )
  );
  X_ZERO   \$4I4029/$1I2653/$1I85/$1I2218  (
    .O(\$4I4029/$1I2653/$1I85/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2653/$1I85/L  (
    .I(\$4I4029/$1I2653/$1I85/$1N2216 ),
    .O(\$4I4029/$1I2653/$1N86 )
  );
  X_ZERO   \$4I4029/$1I2653/$1I88/$1I2218  (
    .O(\$4I4029/$1I2653/$1I88/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2653/$1I88/L  (
    .I(\$4I4029/$1I2653/$1I88/$1N2216 ),
    .O(\$4I4029/$1I2653/$1N87 )
  );
  X_AND2   \$4I4029/$1I2661/$1I31  (
    .I0(\$4I4029/$1N2759 ),
    .I1(\$4I4029/$1I2661/TC ),
    .O(\$4I4029/EXP )
  );
  X_AND4   \$4I4029/$1I2661/$1I28  (
    .I0(\$4I4029/$1I2661/Q6 ),
    .I1(\$4I4029/$1I2661/Q5 ),
    .I2(\$4I4029/$1I2661/Q4 ),
    .I3(\$4I4029/$1I2661/T4 ),
    .O(\$4I4029/$1I2661/T7 )
  );
  X_AND3   \$4I4029/$1I2661/$1I26  (
    .I0(\$4I4029/$1I2661/Q2 ),
    .I1(\$4I4029/$1I2661/Q1 ),
    .I2(\$4I4029/$1I2661/Q0 ),
    .O(\$4I4029/$1I2661/T3 )
  );
  X_AND2   \$4I4029/$1I2661/$1I24  (
    .I0(\$4I4029/$1I2661/Q1 ),
    .I1(\$4I4029/$1I2661/Q0 ),
    .O(\$4I4029/$1I2661/T2 )
  );
  X_AND2   \$4I4029/$1I2661/$1I2  (
    .I0(\$4I4029/$1I2661/Q4 ),
    .I1(\$4I4029/$1I2661/T4 ),
    .O(\$4I4029/$1I2661/T5 )
  );
  X_ONE   \$4I4029/$1I2661/$1I16  (
    .O(\$4I4029/$1I2661/$1N20 )
  );
  X_AND4   \$4I4029/$1I2661/$1I15  (
    .I0(\$4I4029/$1I2661/Q3 ),
    .I1(\$4I4029/$1I2661/Q2 ),
    .I2(\$4I4029/$1I2661/Q1 ),
    .I3(\$4I4029/$1I2661/Q0 ),
    .O(\$4I4029/$1I2661/T4 )
  );
  X_AND3   \$4I4029/$1I2661/$1I11  (
    .I0(\$4I4029/$1I2661/Q5 ),
    .I1(\$4I4029/$1I2661/Q4 ),
    .I2(\$4I4029/$1I2661/T4 ),
    .O(\$4I4029/$1I2661/T6 )
  );
  X_AND5   \$4I4029/$1I2661/$1I1  (
    .I0(\$4I4029/$1I2661/Q7 ),
    .I1(\$4I4029/$1I2661/Q6 ),
    .I2(\$4I4029/$1I2661/Q5 ),
    .I3(\$4I4029/$1I2661/Q4 ),
    .I4(\$4I4029/$1I2661/T4 ),
    .O(\$4I4029/$1I2661/TC )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \$4I4029/$1I2661/$1I43/$1I35  (
    .CE(\$4I4029/$1N2759 ),
    .CLK(CLK),
    .I(\$4I4029/$1I2661/$1I43/MD ),
    .O(\$4I4029/$1I2661/Q0 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \$4I4029/$1I2661/$1I43/$1I32  (
    .I0(\$4I4029/$1I2661/$1N20 ),
    .I1(\$4I4029/$1I2661/Q0 ),
    .O(\$4I4029/$1I2661/$1I43/TQ )
  );
  X_AND2   \$4I4029/$1I2661/$1I43/$1I30/$1I9  (
    .I0(\$4I4029/$1I2661/$1N45 ),
    .I1(\$4I4029/$1I2661/$1N48 ),
    .O(\$4I4029/$1I2661/$1I43/$1I30/M1 )
  );
  X_OR2   \$4I4029/$1I2661/$1I43/$1I30/$1I8  (
    .I0(\$4I4029/$1I2661/$1I43/$1I30/M1 ),
    .I1(\$4I4029/$1I2661/$1I43/$1I30/M0 ),
    .O(\$4I4029/$1I2661/$1I43/MD )
  );
  X_AND2   \$4I4029/$1I2661/$1I43/$1I30/$1I7  (
    .I0(\NlwInverterSignal_$4I4029/$1I2661/$1I43/$1I30/$1I7/I0 ),
    .I1(\$4I4029/$1I2661/$1I43/TQ ),
    .O(\$4I4029/$1I2661/$1I43/$1I30/M0 )
  );
  X_ZERO   \$4I4029/$1I2661/$1I44/$1I2218  (
    .O(\$4I4029/$1I2661/$1I44/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2661/$1I44/L  (
    .I(\$4I4029/$1I2661/$1I44/$1N2216 ),
    .O(\$4I4029/$1I2661/$1N45 )
  );
  X_ZERO   \$4I4029/$1I2661/$1I47/$1I2218  (
    .O(\$4I4029/$1I2661/$1I47/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2661/$1I47/L  (
    .I(\$4I4029/$1I2661/$1I47/$1N2216 ),
    .O(\$4I4029/$1I2661/$1N48 )
  );
  X_ZERO   \$4I4029/$1I2661/$1I49/$1I2218  (
    .O(\$4I4029/$1I2661/$1I49/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2661/$1I49/L  (
    .I(\$4I4029/$1I2661/$1I49/$1N2216 ),
    .O(\$4I4029/$1I2661/$1N50 )
  );
  X_ZERO   \$4I4029/$1I2661/$1I52/$1I2218  (
    .O(\$4I4029/$1I2661/$1I52/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2661/$1I52/L  (
    .I(\$4I4029/$1I2661/$1I52/$1N2216 ),
    .O(\$4I4029/$1I2661/$1N51 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \$4I4029/$1I2661/$1I53/$1I35  (
    .CE(\$4I4029/$1N2759 ),
    .CLK(CLK),
    .I(\$4I4029/$1I2661/$1I53/MD ),
    .O(\$4I4029/$1I2661/Q1 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \$4I4029/$1I2661/$1I53/$1I32  (
    .I0(\$4I4029/$1I2661/Q0 ),
    .I1(\$4I4029/$1I2661/Q1 ),
    .O(\$4I4029/$1I2661/$1I53/TQ )
  );
  X_AND2   \$4I4029/$1I2661/$1I53/$1I30/$1I9  (
    .I0(\$4I4029/$1I2661/$1N50 ),
    .I1(\$4I4029/$1I2661/$1N51 ),
    .O(\$4I4029/$1I2661/$1I53/$1I30/M1 )
  );
  X_OR2   \$4I4029/$1I2661/$1I53/$1I30/$1I8  (
    .I0(\$4I4029/$1I2661/$1I53/$1I30/M1 ),
    .I1(\$4I4029/$1I2661/$1I53/$1I30/M0 ),
    .O(\$4I4029/$1I2661/$1I53/MD )
  );
  X_AND2   \$4I4029/$1I2661/$1I53/$1I30/$1I7  (
    .I0(\NlwInverterSignal_$4I4029/$1I2661/$1I53/$1I30/$1I7/I0 ),
    .I1(\$4I4029/$1I2661/$1I53/TQ ),
    .O(\$4I4029/$1I2661/$1I53/$1I30/M0 )
  );
  X_ZERO   \$4I4029/$1I2661/$1I54/$1I2218  (
    .O(\$4I4029/$1I2661/$1I54/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2661/$1I54/L  (
    .I(\$4I4029/$1I2661/$1I54/$1N2216 ),
    .O(\$4I4029/$1I2661/$1N55 )
  );
  X_ZERO   \$4I4029/$1I2661/$1I57/$1I2218  (
    .O(\$4I4029/$1I2661/$1I57/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2661/$1I57/L  (
    .I(\$4I4029/$1I2661/$1I57/$1N2216 ),
    .O(\$4I4029/$1I2661/$1N56 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \$4I4029/$1I2661/$1I58/$1I35  (
    .CE(\$4I4029/$1N2759 ),
    .CLK(CLK),
    .I(\$4I4029/$1I2661/$1I58/MD ),
    .O(\$4I4029/$1I2661/Q2 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \$4I4029/$1I2661/$1I58/$1I32  (
    .I0(\$4I4029/$1I2661/T2 ),
    .I1(\$4I4029/$1I2661/Q2 ),
    .O(\$4I4029/$1I2661/$1I58/TQ )
  );
  X_AND2   \$4I4029/$1I2661/$1I58/$1I30/$1I9  (
    .I0(\$4I4029/$1I2661/$1N55 ),
    .I1(\$4I4029/$1I2661/$1N56 ),
    .O(\$4I4029/$1I2661/$1I58/$1I30/M1 )
  );
  X_OR2   \$4I4029/$1I2661/$1I58/$1I30/$1I8  (
    .I0(\$4I4029/$1I2661/$1I58/$1I30/M1 ),
    .I1(\$4I4029/$1I2661/$1I58/$1I30/M0 ),
    .O(\$4I4029/$1I2661/$1I58/MD )
  );
  X_AND2   \$4I4029/$1I2661/$1I58/$1I30/$1I7  (
    .I0(\NlwInverterSignal_$4I4029/$1I2661/$1I58/$1I30/$1I7/I0 ),
    .I1(\$4I4029/$1I2661/$1I58/TQ ),
    .O(\$4I4029/$1I2661/$1I58/$1I30/M0 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \$4I4029/$1I2661/$1I59/$1I35  (
    .CE(\$4I4029/$1N2759 ),
    .CLK(CLK),
    .I(\$4I4029/$1I2661/$1I59/MD ),
    .O(\$4I4029/$1I2661/Q3 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \$4I4029/$1I2661/$1I59/$1I32  (
    .I0(\$4I4029/$1I2661/T3 ),
    .I1(\$4I4029/$1I2661/Q3 ),
    .O(\$4I4029/$1I2661/$1I59/TQ )
  );
  X_AND2   \$4I4029/$1I2661/$1I59/$1I30/$1I9  (
    .I0(\$4I4029/$1I2661/$1N62 ),
    .I1(\$4I4029/$1I2661/$1N61 ),
    .O(\$4I4029/$1I2661/$1I59/$1I30/M1 )
  );
  X_OR2   \$4I4029/$1I2661/$1I59/$1I30/$1I8  (
    .I0(\$4I4029/$1I2661/$1I59/$1I30/M1 ),
    .I1(\$4I4029/$1I2661/$1I59/$1I30/M0 ),
    .O(\$4I4029/$1I2661/$1I59/MD )
  );
  X_AND2   \$4I4029/$1I2661/$1I59/$1I30/$1I7  (
    .I0(\NlwInverterSignal_$4I4029/$1I2661/$1I59/$1I30/$1I7/I0 ),
    .I1(\$4I4029/$1I2661/$1I59/TQ ),
    .O(\$4I4029/$1I2661/$1I59/$1I30/M0 )
  );
  X_ZERO   \$4I4029/$1I2661/$1I60/$1I2218  (
    .O(\$4I4029/$1I2661/$1I60/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2661/$1I60/L  (
    .I(\$4I4029/$1I2661/$1I60/$1N2216 ),
    .O(\$4I4029/$1I2661/$1N61 )
  );
  X_ZERO   \$4I4029/$1I2661/$1I63/$1I2218  (
    .O(\$4I4029/$1I2661/$1I63/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2661/$1I63/L  (
    .I(\$4I4029/$1I2661/$1I63/$1N2216 ),
    .O(\$4I4029/$1I2661/$1N62 )
  );
  X_ZERO   \$4I4029/$1I2661/$1I64/$1I2218  (
    .O(\$4I4029/$1I2661/$1I64/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2661/$1I64/L  (
    .I(\$4I4029/$1I2661/$1I64/$1N2216 ),
    .O(\$4I4029/$1I2661/$1N65 )
  );
  X_ZERO   \$4I4029/$1I2661/$1I67/$1I2218  (
    .O(\$4I4029/$1I2661/$1I67/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2661/$1I67/L  (
    .I(\$4I4029/$1I2661/$1I67/$1N2216 ),
    .O(\$4I4029/$1I2661/$1N66 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \$4I4029/$1I2661/$1I68/$1I35  (
    .CE(\$4I4029/$1N2759 ),
    .CLK(CLK),
    .I(\$4I4029/$1I2661/$1I68/MD ),
    .O(\$4I4029/$1I2661/Q4 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \$4I4029/$1I2661/$1I68/$1I32  (
    .I0(\$4I4029/$1I2661/T4 ),
    .I1(\$4I4029/$1I2661/Q4 ),
    .O(\$4I4029/$1I2661/$1I68/TQ )
  );
  X_AND2   \$4I4029/$1I2661/$1I68/$1I30/$1I9  (
    .I0(\$4I4029/$1I2661/$1N65 ),
    .I1(\$4I4029/$1I2661/$1N66 ),
    .O(\$4I4029/$1I2661/$1I68/$1I30/M1 )
  );
  X_OR2   \$4I4029/$1I2661/$1I68/$1I30/$1I8  (
    .I0(\$4I4029/$1I2661/$1I68/$1I30/M1 ),
    .I1(\$4I4029/$1I2661/$1I68/$1I30/M0 ),
    .O(\$4I4029/$1I2661/$1I68/MD )
  );
  X_AND2   \$4I4029/$1I2661/$1I68/$1I30/$1I7  (
    .I0(\NlwInverterSignal_$4I4029/$1I2661/$1I68/$1I30/$1I7/I0 ),
    .I1(\$4I4029/$1I2661/$1I68/TQ ),
    .O(\$4I4029/$1I2661/$1I68/$1I30/M0 )
  );
  X_ZERO   \$4I4029/$1I2661/$1I69/$1I2218  (
    .O(\$4I4029/$1I2661/$1I69/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2661/$1I69/L  (
    .I(\$4I4029/$1I2661/$1I69/$1N2216 ),
    .O(\$4I4029/$1I2661/$1N70 )
  );
  X_ZERO   \$4I4029/$1I2661/$1I72/$1I2218  (
    .O(\$4I4029/$1I2661/$1I72/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2661/$1I72/L  (
    .I(\$4I4029/$1I2661/$1I72/$1N2216 ),
    .O(\$4I4029/$1I2661/$1N71 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \$4I4029/$1I2661/$1I73/$1I35  (
    .CE(\$4I4029/$1N2759 ),
    .CLK(CLK),
    .I(\$4I4029/$1I2661/$1I73/MD ),
    .O(\$4I4029/$1I2661/Q5 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \$4I4029/$1I2661/$1I73/$1I32  (
    .I0(\$4I4029/$1I2661/T5 ),
    .I1(\$4I4029/$1I2661/Q5 ),
    .O(\$4I4029/$1I2661/$1I73/TQ )
  );
  X_AND2   \$4I4029/$1I2661/$1I73/$1I30/$1I9  (
    .I0(\$4I4029/$1I2661/$1N70 ),
    .I1(\$4I4029/$1I2661/$1N71 ),
    .O(\$4I4029/$1I2661/$1I73/$1I30/M1 )
  );
  X_OR2   \$4I4029/$1I2661/$1I73/$1I30/$1I8  (
    .I0(\$4I4029/$1I2661/$1I73/$1I30/M1 ),
    .I1(\$4I4029/$1I2661/$1I73/$1I30/M0 ),
    .O(\$4I4029/$1I2661/$1I73/MD )
  );
  X_AND2   \$4I4029/$1I2661/$1I73/$1I30/$1I7  (
    .I0(\NlwInverterSignal_$4I4029/$1I2661/$1I73/$1I30/$1I7/I0 ),
    .I1(\$4I4029/$1I2661/$1I73/TQ ),
    .O(\$4I4029/$1I2661/$1I73/$1I30/M0 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \$4I4029/$1I2661/$1I79/$1I35  (
    .CE(\$4I4029/$1N2759 ),
    .CLK(CLK),
    .I(\$4I4029/$1I2661/$1I79/MD ),
    .O(\$4I4029/$1I2661/Q6 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \$4I4029/$1I2661/$1I79/$1I32  (
    .I0(\$4I4029/$1I2661/T6 ),
    .I1(\$4I4029/$1I2661/Q6 ),
    .O(\$4I4029/$1I2661/$1I79/TQ )
  );
  X_AND2   \$4I4029/$1I2661/$1I79/$1I30/$1I9  (
    .I0(\$4I4029/$1I2661/$1N82 ),
    .I1(\$4I4029/$1I2661/$1N81 ),
    .O(\$4I4029/$1I2661/$1I79/$1I30/M1 )
  );
  X_OR2   \$4I4029/$1I2661/$1I79/$1I30/$1I8  (
    .I0(\$4I4029/$1I2661/$1I79/$1I30/M1 ),
    .I1(\$4I4029/$1I2661/$1I79/$1I30/M0 ),
    .O(\$4I4029/$1I2661/$1I79/MD )
  );
  X_AND2   \$4I4029/$1I2661/$1I79/$1I30/$1I7  (
    .I0(\NlwInverterSignal_$4I4029/$1I2661/$1I79/$1I30/$1I7/I0 ),
    .I1(\$4I4029/$1I2661/$1I79/TQ ),
    .O(\$4I4029/$1I2661/$1I79/$1I30/M0 )
  );
  X_ZERO   \$4I4029/$1I2661/$1I80/$1I2218  (
    .O(\$4I4029/$1I2661/$1I80/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2661/$1I80/L  (
    .I(\$4I4029/$1I2661/$1I80/$1N2216 ),
    .O(\$4I4029/$1I2661/$1N81 )
  );
  X_ZERO   \$4I4029/$1I2661/$1I83/$1I2218  (
    .O(\$4I4029/$1I2661/$1I83/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2661/$1I83/L  (
    .I(\$4I4029/$1I2661/$1I83/$1N2216 ),
    .O(\$4I4029/$1I2661/$1N82 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \$4I4029/$1I2661/$1I84/$1I35  (
    .CE(\$4I4029/$1N2759 ),
    .CLK(CLK),
    .I(\$4I4029/$1I2661/$1I84/MD ),
    .O(\$4I4029/$1I2661/Q7 ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_XOR2   \$4I4029/$1I2661/$1I84/$1I32  (
    .I0(\$4I4029/$1I2661/T7 ),
    .I1(\$4I4029/$1I2661/Q7 ),
    .O(\$4I4029/$1I2661/$1I84/TQ )
  );
  X_AND2   \$4I4029/$1I2661/$1I84/$1I30/$1I9  (
    .I0(\$4I4029/$1I2661/$1N87 ),
    .I1(\$4I4029/$1I2661/$1N86 ),
    .O(\$4I4029/$1I2661/$1I84/$1I30/M1 )
  );
  X_OR2   \$4I4029/$1I2661/$1I84/$1I30/$1I8  (
    .I0(\$4I4029/$1I2661/$1I84/$1I30/M1 ),
    .I1(\$4I4029/$1I2661/$1I84/$1I30/M0 ),
    .O(\$4I4029/$1I2661/$1I84/MD )
  );
  X_AND2   \$4I4029/$1I2661/$1I84/$1I30/$1I7  (
    .I0(\NlwInverterSignal_$4I4029/$1I2661/$1I84/$1I30/$1I7/I0 ),
    .I1(\$4I4029/$1I2661/$1I84/TQ ),
    .O(\$4I4029/$1I2661/$1I84/$1I30/M0 )
  );
  X_ZERO   \$4I4029/$1I2661/$1I85/$1I2218  (
    .O(\$4I4029/$1I2661/$1I85/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2661/$1I85/L  (
    .I(\$4I4029/$1I2661/$1I85/$1N2216 ),
    .O(\$4I4029/$1I2661/$1N86 )
  );
  X_ZERO   \$4I4029/$1I2661/$1I88/$1I2218  (
    .O(\$4I4029/$1I2661/$1I88/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2661/$1I88/L  (
    .I(\$4I4029/$1I2661/$1I88/$1N2216 ),
    .O(\$4I4029/$1I2661/$1N87 )
  );
  X_ONE   \$4I4029/$1I2730/$1I2220  (
    .O(\$4I4029/$1I2730/$1N2216 )
  );
  X_BUF   \$4I4029/$1I2730/H  (
    .I(\$4I4029/$1I2730/$1N2216 ),
    .O(\$4I4029/ONE )
  );
  X_ZERO   \$4I4076/$1I2218  (
    .O(\$4I4076/$1N2216 )
  );
  X_BUF   \$4I4076/L  (
    .I(\$4I4076/$1N2216 ),
    .O(SET6)
  );
  X_ZERO   \$4I4095/$1I2218  (
    .O(\$4I4095/$1N2216 )
  );
  X_BUF   \$4I4095/L  (
    .I(\$4I4095/$1N2216 ),
    .O(SET9)
  );
  X_ZERO   \$4I4096/$1I2218  (
    .O(\$4I4096/$1N2216 )
  );
  X_BUF   \$4I4096/L  (
    .I(\$4I4096/$1N2216 ),
    .O(SET7)
  );
  X_ZERO   \$4I4097/$1I2218  (
    .O(\$4I4097/$1N2216 )
  );
  X_BUF   \$4I4097/L  (
    .I(\$4I4097/$1N2216 ),
    .O(SET5)
  );
  X_ZERO   \$4I4098/$1I2218  (
    .O(\$4I4098/$1N2216 )
  );
  X_BUF   \$4I4098/L  (
    .I(\$4I4098/$1N2216 ),
    .O(SET4)
  );
  X_ZERO   \$4I4099/$1I2218  (
    .O(\$4I4099/$1N2216 )
  );
  X_BUF   \$4I4099/L  (
    .I(\$4I4099/$1N2216 ),
    .O(SET3)
  );
  X_ZERO   \$4I4100/$1I2218  (
    .O(\$4I4100/$1N2216 )
  );
  X_BUF   \$4I4100/L  (
    .I(\$4I4100/$1N2216 ),
    .O(SET2)
  );
  X_ZERO   \$4I4101/$1I2218  (
    .O(\$4I4101/$1N2216 )
  );
  X_BUF   \$4I4101/L  (
    .I(\$4I4101/$1N2216 ),
    .O(SET1)
  );
  X_ZERO   \$4I4102/$1I2218  (
    .O(\$4I4102/$1N2216 )
  );
  X_BUF   \$4I4102/L  (
    .I(\$4I4102/$1N2216 ),
    .O(SET10)
  );
  X_ZERO   \$4I4103/$1I2218  (
    .O(\$4I4103/$1N2216 )
  );
  X_BUF   \$4I4103/L  (
    .I(\$4I4103/$1N2216 ),
    .O(SET0)
  );
  X_TRI   \E/UPPER/T0  (
    .I(AD16),
    .O(ADIO16),
    .CTL(\NlwInverterSignal_E/UPPER/T0/T )
  );
  X_TRI   \E/UPPER/T1  (
    .I(AD17),
    .O(ADIO17),
    .CTL(\NlwInverterSignal_E/UPPER/T1/T )
  );
  X_TRI   \E/UPPER/T2  (
    .I(AD18),
    .O(ADIO18),
    .CTL(\NlwInverterSignal_E/UPPER/T2/T )
  );
  X_TRI   \E/UPPER/T3  (
    .I(AD19),
    .O(ADIO19),
    .CTL(\NlwInverterSignal_E/UPPER/T3/T )
  );
  X_TRI   \E/UPPER/T4  (
    .I(AD20),
    .O(ADIO20),
    .CTL(\NlwInverterSignal_E/UPPER/T4/T )
  );
  X_TRI   \E/UPPER/T5  (
    .I(AD21),
    .O(ADIO21),
    .CTL(\NlwInverterSignal_E/UPPER/T5/T )
  );
  X_TRI   \E/UPPER/T6  (
    .I(AD22),
    .O(ADIO22),
    .CTL(\NlwInverterSignal_E/UPPER/T6/T )
  );
  X_TRI   \E/UPPER/T7  (
    .I(AD23),
    .O(ADIO23),
    .CTL(\NlwInverterSignal_E/UPPER/T7/T )
  );
  X_TRI   \E/UPPER/T8  (
    .I(AD24),
    .O(ADIO24),
    .CTL(\NlwInverterSignal_E/UPPER/T8/T )
  );
  X_TRI   \E/UPPER/T9  (
    .I(AD25),
    .O(ADIO25),
    .CTL(\NlwInverterSignal_E/UPPER/T9/T )
  );
  X_TRI   \E/UPPER/T10  (
    .I(AD26),
    .O(ADIO26),
    .CTL(\NlwInverterSignal_E/UPPER/T10/T )
  );
  X_TRI   \E/UPPER/T11  (
    .I(AD27),
    .O(ADIO27),
    .CTL(\NlwInverterSignal_E/UPPER/T11/T )
  );
  X_TRI   \E/UPPER/T12  (
    .I(AD28),
    .O(ADIO28),
    .CTL(\NlwInverterSignal_E/UPPER/T12/T )
  );
  X_TRI   \E/UPPER/T13  (
    .I(AD29),
    .O(ADIO29),
    .CTL(\NlwInverterSignal_E/UPPER/T13/T )
  );
  X_TRI   \E/UPPER/T14  (
    .I(AD30),
    .O(ADIO30),
    .CTL(\NlwInverterSignal_E/UPPER/T14/T )
  );
  X_TRI   \E/UPPER/T15  (
    .I(AD31),
    .O(ADIO31),
    .CTL(\NlwInverterSignal_E/UPPER/T15/T )
  );
  X_TRI   \E/LOWER/T0  (
    .I(AD0),
    .O(ADIO0),
    .CTL(\NlwInverterSignal_E/LOWER/T0/T )
  );
  X_TRI   \E/LOWER/T1  (
    .I(AD1),
    .O(ADIO1),
    .CTL(\NlwInverterSignal_E/LOWER/T1/T )
  );
  X_TRI   \E/LOWER/T2  (
    .I(AD2),
    .O(ADIO2),
    .CTL(\NlwInverterSignal_E/LOWER/T2/T )
  );
  X_TRI   \E/LOWER/T3  (
    .I(AD3),
    .O(ADIO3),
    .CTL(\NlwInverterSignal_E/LOWER/T3/T )
  );
  X_TRI   \E/LOWER/T4  (
    .I(AD4),
    .O(ADIO4),
    .CTL(\NlwInverterSignal_E/LOWER/T4/T )
  );
  X_TRI   \E/LOWER/T5  (
    .I(AD5),
    .O(ADIO5),
    .CTL(\NlwInverterSignal_E/LOWER/T5/T )
  );
  X_TRI   \E/LOWER/T6  (
    .I(AD6),
    .O(ADIO6),
    .CTL(\NlwInverterSignal_E/LOWER/T6/T )
  );
  X_TRI   \E/LOWER/T7  (
    .I(AD7),
    .O(ADIO7),
    .CTL(\NlwInverterSignal_E/LOWER/T7/T )
  );
  X_TRI   \E/LOWER/T8  (
    .I(AD8),
    .O(ADIO8),
    .CTL(\NlwInverterSignal_E/LOWER/T8/T )
  );
  X_TRI   \E/LOWER/T9  (
    .I(AD9),
    .O(ADIO9),
    .CTL(\NlwInverterSignal_E/LOWER/T9/T )
  );
  X_TRI   \E/LOWER/T10  (
    .I(AD10),
    .O(ADIO10),
    .CTL(\NlwInverterSignal_E/LOWER/T10/T )
  );
  X_TRI   \E/LOWER/T11  (
    .I(AD11),
    .O(ADIO11),
    .CTL(\NlwInverterSignal_E/LOWER/T11/T )
  );
  X_TRI   \E/LOWER/T12  (
    .I(AD12),
    .O(ADIO12),
    .CTL(\NlwInverterSignal_E/LOWER/T12/T )
  );
  X_TRI   \E/LOWER/T13  (
    .I(AD13),
    .O(ADIO13),
    .CTL(\NlwInverterSignal_E/LOWER/T13/T )
  );
  X_TRI   \E/LOWER/T14  (
    .I(AD14),
    .O(ADIO14),
    .CTL(\NlwInverterSignal_E/LOWER/T14/T )
  );
  X_TRI   \E/LOWER/T15  (
    .I(AD15),
    .O(ADIO15),
    .CTL(\NlwInverterSignal_E/LOWER/T15/T )
  );
  X_TRI   \E64/UPPER/T0  (
    .I(AD48),
    .O(ADIO48),
    .CTL(\NlwInverterSignal_E64/UPPER/T0/T )
  );
  X_TRI   \E64/UPPER/T1  (
    .I(AD49),
    .O(ADIO49),
    .CTL(\NlwInverterSignal_E64/UPPER/T1/T )
  );
  X_TRI   \E64/UPPER/T2  (
    .I(AD50),
    .O(ADIO50),
    .CTL(\NlwInverterSignal_E64/UPPER/T2/T )
  );
  X_TRI   \E64/UPPER/T3  (
    .I(AD51),
    .O(ADIO51),
    .CTL(\NlwInverterSignal_E64/UPPER/T3/T )
  );
  X_TRI   \E64/UPPER/T4  (
    .I(AD52),
    .O(ADIO52),
    .CTL(\NlwInverterSignal_E64/UPPER/T4/T )
  );
  X_TRI   \E64/UPPER/T5  (
    .I(AD53),
    .O(ADIO53),
    .CTL(\NlwInverterSignal_E64/UPPER/T5/T )
  );
  X_TRI   \E64/UPPER/T6  (
    .I(AD54),
    .O(ADIO54),
    .CTL(\NlwInverterSignal_E64/UPPER/T6/T )
  );
  X_TRI   \E64/UPPER/T7  (
    .I(AD55),
    .O(ADIO55),
    .CTL(\NlwInverterSignal_E64/UPPER/T7/T )
  );
  X_TRI   \E64/UPPER/T8  (
    .I(AD56),
    .O(ADIO56),
    .CTL(\NlwInverterSignal_E64/UPPER/T8/T )
  );
  X_TRI   \E64/UPPER/T9  (
    .I(AD57),
    .O(ADIO57),
    .CTL(\NlwInverterSignal_E64/UPPER/T9/T )
  );
  X_TRI   \E64/UPPER/T10  (
    .I(AD58),
    .O(ADIO58),
    .CTL(\NlwInverterSignal_E64/UPPER/T10/T )
  );
  X_TRI   \E64/UPPER/T11  (
    .I(AD59),
    .O(ADIO59),
    .CTL(\NlwInverterSignal_E64/UPPER/T11/T )
  );
  X_TRI   \E64/UPPER/T12  (
    .I(AD60),
    .O(ADIO60),
    .CTL(\NlwInverterSignal_E64/UPPER/T12/T )
  );
  X_TRI   \E64/UPPER/T13  (
    .I(AD61),
    .O(ADIO61),
    .CTL(\NlwInverterSignal_E64/UPPER/T13/T )
  );
  X_TRI   \E64/UPPER/T14  (
    .I(AD62),
    .O(ADIO62),
    .CTL(\NlwInverterSignal_E64/UPPER/T14/T )
  );
  X_TRI   \E64/UPPER/T15  (
    .I(AD63),
    .O(ADIO63),
    .CTL(\NlwInverterSignal_E64/UPPER/T15/T )
  );
  X_TRI   \E64/LOWER/T0  (
    .I(AD32),
    .O(ADIO32),
    .CTL(\NlwInverterSignal_E64/LOWER/T0/T )
  );
  X_TRI   \E64/LOWER/T1  (
    .I(AD33),
    .O(ADIO33),
    .CTL(\NlwInverterSignal_E64/LOWER/T1/T )
  );
  X_TRI   \E64/LOWER/T2  (
    .I(AD34),
    .O(ADIO34),
    .CTL(\NlwInverterSignal_E64/LOWER/T2/T )
  );
  X_TRI   \E64/LOWER/T3  (
    .I(AD35),
    .O(ADIO35),
    .CTL(\NlwInverterSignal_E64/LOWER/T3/T )
  );
  X_TRI   \E64/LOWER/T4  (
    .I(AD36),
    .O(ADIO36),
    .CTL(\NlwInverterSignal_E64/LOWER/T4/T )
  );
  X_TRI   \E64/LOWER/T5  (
    .I(AD37),
    .O(ADIO37),
    .CTL(\NlwInverterSignal_E64/LOWER/T5/T )
  );
  X_TRI   \E64/LOWER/T6  (
    .I(AD38),
    .O(ADIO38),
    .CTL(\NlwInverterSignal_E64/LOWER/T6/T )
  );
  X_TRI   \E64/LOWER/T7  (
    .I(AD39),
    .O(ADIO39),
    .CTL(\NlwInverterSignal_E64/LOWER/T7/T )
  );
  X_TRI   \E64/LOWER/T8  (
    .I(AD40),
    .O(ADIO40),
    .CTL(\NlwInverterSignal_E64/LOWER/T8/T )
  );
  X_TRI   \E64/LOWER/T9  (
    .I(AD41),
    .O(ADIO41),
    .CTL(\NlwInverterSignal_E64/LOWER/T9/T )
  );
  X_TRI   \E64/LOWER/T10  (
    .I(AD42),
    .O(ADIO42),
    .CTL(\NlwInverterSignal_E64/LOWER/T10/T )
  );
  X_TRI   \E64/LOWER/T11  (
    .I(AD43),
    .O(ADIO43),
    .CTL(\NlwInverterSignal_E64/LOWER/T11/T )
  );
  X_TRI   \E64/LOWER/T12  (
    .I(AD44),
    .O(ADIO44),
    .CTL(\NlwInverterSignal_E64/LOWER/T12/T )
  );
  X_TRI   \E64/LOWER/T13  (
    .I(AD45),
    .O(ADIO45),
    .CTL(\NlwInverterSignal_E64/LOWER/T13/T )
  );
  X_TRI   \E64/LOWER/T14  (
    .I(AD46),
    .O(ADIO46),
    .CTL(\NlwInverterSignal_E64/LOWER/T14/T )
  );
  X_TRI   \E64/LOWER/T15  (
    .I(AD47),
    .O(ADIO47),
    .CTL(\NlwInverterSignal_E64/LOWER/T15/T )
  );
  X_AND2   \OEADI/$1I4041  (
    .I0(\NlwInverterSignal_OEADI/$1I4041/I0 ),
    .I1(S_WRDN_DUP),
    .O(\OEADI/$1N4030 )
  );
  X_AND2   \OEADI/$1I4040  (
    .I0(\NlwInverterSignal_OEADI/$1I4040/I0 ),
    .I1(IDLE_DUP),
    .O(\OEADI/$1N4036 )
  );
  X_MUX2   \OEADI/$1I4037  (
    .IA(\OEADI/OAI64_0 ),
    .IB(\OEADI/OAI64_1 ),
    .O(OE_ADI64),
    .SEL(I_IDLE_INT)
  );
  X_AND4   \OEADI/$1I4031  (
    .I0(\NlwInverterSignal_OEADI/$1I4031/I0 ),
    .I1(\NlwInverterSignal_OEADI/$1I4031/I1 ),
    .I2(\NlwInverterSignal_OEADI/$1I4031/I2 ),
    .I3(M_DATA_INT),
    .O(\NlwInverterSignal_OEADI/$1I4031/O )
  );
  X_OR2   \OEADI/$1I4029  (
    .I0(\OEADI/$1N4036 ),
    .I1(\OEADI/$1N4030 ),
    .O(\OEADI/$1N4042 )
  );
  X_AND2   \OEADI/$1I4028  (
    .I0(\NlwInverterSignal_OEADI/$1I4028/I0 ),
    .I1(\OEADI/$1N4042 ),
    .O(\NlwInverterSignal_OEADI/$1I4028/O )
  );
  X_OR3   \OEADI/$1I3995  (
    .I0(\OEADI/M_DATAQ ),
    .I1(OLDKEEPOUT),
    .I2(ADDR_BE),
    .O(\OEADI/MIDDLE )
  );
  X_AND2   \OEADI/$1I3984  (
    .I0(\NlwInverterSignal_OEADI/$1I3984/I0 ),
    .I1(\OEADI/$1N3986 ),
    .O(\NlwInverterSignal_OEADI/$1I3984/O )
  );
  X_OR2   \OEADI/$1I3983  (
    .I0(\OEADI/$1N3857 ),
    .I1(\OEADI/$1N3855 ),
    .O(\OEADI/$1N3986 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \OEADI/CSQ_FF  (
    .CE(VCC),
    .CLK(CLK),
    .I(CFG_SELF),
    .O(\OEADI/CFG_SELFQ ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_AND4   \OEADI/$1I3954  (
    .I0(\NlwInverterSignal_OEADI/$1I3954/I0 ),
    .I1(\NlwInverterSignal_OEADI/$1I3954/I1 ),
    .I2(\NlwInverterSignal_OEADI/$1I3954/I2 ),
    .I3(M_DATA_INT),
    .O(\NlwInverterSignal_OEADI/$1I3954/O )
  );
  X_MUX2   \OEADI/$1I3951  (
    .IA(\OEADI/OAI32_0 ),
    .IB(\OEADI/OAI32_1 ),
    .O(OE_ADI),
    .SEL(I_IDLE_INT)
  );
  X_AND2   \OEADI/$1I3864  (
    .I0(\NlwInverterSignal_OEADI/$1I3864/I0 ),
    .I1(IDLE_DUP),
    .O(\OEADI/$1N3857 )
  );
  X_AND2   \OEADI/$1I3860  (
    .I0(\NlwInverterSignal_OEADI/$1I3860/I0 ),
    .I1(S_WRDN_DUP),
    .O(\OEADI/$1N3855 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \OEADI/MDQ_FF  (
    .CE(VCC),
    .CLK(CLK),
    .I(M_DATA_INT),
    .O(\OEADI/M_DATAQ ),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_BUF   \OEADI/$1I4047/NC  (
    .I(DR_BUS_INT),
    .O(\NLW_OEADI/$1I4047/NC_O_UNCONNECTED )
  );
  X_AND2   \$5I3771/$1I9  (
    .I0(\$5N3772 ),
    .I1(CFG111),
    .O(\$5I3771/M1 )
  );
  X_OR2   \$5I3771/$1I8  (
    .I0(\$5I3771/M1 ),
    .I1(\$5I3771/M0 ),
    .O(OLDKEEPOUT)
  );
  X_AND2   \$5I3771/$1I7  (
    .I0(\NlwInverterSignal_$5I3771/$1I7/I0 ),
    .I1(KEEPOUT),
    .O(\$5I3771/M0 )
  );
  X_ZERO   \$5I3778/$1I2218  (
    .O(\$5I3778/$1N2216 )
  );
  X_BUF   \$5I3778/L  (
    .I(\$5I3778/$1N2216 ),
    .O(\$5N3772 )
  );
  X_AND2   \$5I3781/$1I9  (
    .I0(KEEPOUT),
    .I1(CFG111),
    .O(\$5I3781/M1 )
  );
  X_OR2   \$5I3781/$1I8  (
    .I0(\$5I3781/M1 ),
    .I1(\$5I3781/M0 ),
    .O(MIKELOVEJOY)
  );
  X_AND2   \$5I3781/$1I7  (
    .I0(\NlwInverterSignal_$5I3781/$1I7/I0 ),
    .I1(\$5N3783 ),
    .O(\$5I3781/M0 )
  );
  X_ZERO   \$5I3782/$1I2218  (
    .O(\$5I3782/$1N2216 )
  );
  X_BUF   \$5I3782/L  (
    .I(\$5I3782/$1N2216 ),
    .O(\$5N3783 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PAR64/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PAR_CE),
    .CLK(CLK),
    .I(NS_PAR64),
    .O(PAR64_O),
    .RST(GND)
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PAR/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PAR_CE),
    .CLK(CLK),
    .I(NS_PAR),
    .O(PAR_O),
    .RST(GND)
  );
  X_BUF   \$6I1087/NC  (
    .I(IDSEL_O),
    .O(\NLW_$6I1087/NC_O_UNCONNECTED )
  );
  X_BUF   \$6I1090/NC  (
    .I(SERR_O),
    .O(\NLW_$6I1090/NC_O_UNCONNECTED )
  );
  X_BUF   \DEVSEL/$1I2284  (
    .I(DEVSEL_I),
    .O(\DEVSEL/D1_9541 )
  );
  X_BUF   \DEVSEL/$1I2282  (
    .I(\DEVSEL/D1_9541 ),
    .O(\DEVSEL/D2_9539 )
  );
  X_BUF   \DEVSEL/$1I2281  (
    .I(\DEVSEL/D2_9539 ),
    .O(\DEVSEL/D3_9540 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \DEVSEL/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(DEVSEL_CE),
    .CLK(CLK),
    .I(\NS_DEVSEL- ),
    .O(DEVSEL_O),
    .RST(GND)
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \DEVSEL/IFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(\DEVSEL/$1N2275 ),
    .CLK(CLK),
    .I(\DEVSEL/IN ),
    .O(\DEVSEL- ),
    .RST(GND)
  );
  X_ONE   \DEVSEL/$1I2276/$1I2220  (
    .O(\DEVSEL/$1I2276/$1N2216 )
  );
  X_BUF   \DEVSEL/$1I2276/H  (
    .I(\DEVSEL/$1I2276/$1N2216 ),
    .O(\DEVSEL/$1N2275 )
  );
  X_ONE   \DEVSEL/$1I2306/$1I2220  (
    .O(\DEVSEL/$1I2306/$1N2216 )
  );
  X_BUF   \DEVSEL/$1I2306/H  (
    .I(\DEVSEL/$1I2306/$1N2216 ),
    .O(\DEVSEL/$1N2307 )
  );
  X_MUX2   \DEVSEL/$1I2310/O  (
    .IA(\DEVSEL/$1I2310/M01 ),
    .IB(\DEVSEL/$1I2310/M23 ),
    .O(\DEVSEL/IN ),
    .SEL(CFG248)
  );
  X_OR2   \DEVSEL/$1I2310/M01/$1I38  (
    .I0(\DEVSEL/$1I2310/M01/M1 ),
    .I1(\DEVSEL/$1I2310/M01/M0 ),
    .O(\DEVSEL/$1I2310/M01 )
  );
  X_AND3   \DEVSEL/$1I2310/M01/$1I31  (
    .I0(\NlwInverterSignal_DEVSEL/$1I2310/M01/$1I31/I0 ),
    .I1(\DEVSEL/$1N2307 ),
    .I2(DEVSEL_I),
    .O(\DEVSEL/$1I2310/M01/M0 )
  );
  X_AND3   \DEVSEL/$1I2310/M01/$1I30  (
    .I0(\DEVSEL/D1_9541 ),
    .I1(\DEVSEL/$1N2307 ),
    .I2(CFG247),
    .O(\DEVSEL/$1I2310/M01/M1 )
  );
  X_OR2   \DEVSEL/$1I2310/M23/$1I38  (
    .I0(\DEVSEL/$1I2310/M23/M1 ),
    .I1(\DEVSEL/$1I2310/M23/M0 ),
    .O(\DEVSEL/$1I2310/M23 )
  );
  X_AND3   \DEVSEL/$1I2310/M23/$1I31  (
    .I0(\NlwInverterSignal_DEVSEL/$1I2310/M23/$1I31/I0 ),
    .I1(\DEVSEL/$1N2307 ),
    .I2(\DEVSEL/D2_9539 ),
    .O(\DEVSEL/$1I2310/M23/M0 )
  );
  X_AND3   \DEVSEL/$1I2310/M23/$1I30  (
    .I0(\DEVSEL/D3_9540 ),
    .I1(\DEVSEL/$1N2307 ),
    .I2(CFG247),
    .O(\DEVSEL/$1I2310/M23/M1 )
  );
  X_BUF   \ACK64/$1I2284  (
    .I(ACK64_I),
    .O(\ACK64/D1_9585 )
  );
  X_BUF   \ACK64/$1I2282  (
    .I(\ACK64/D1_9585 ),
    .O(\ACK64/D2_9583 )
  );
  X_BUF   \ACK64/$1I2281  (
    .I(\ACK64/D2_9583 ),
    .O(\ACK64/D3_9584 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \ACK64/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(ACK64_CE),
    .CLK(CLK),
    .I(\NS_ACK64- ),
    .O(ACK64_O),
    .RST(GND)
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \ACK64/IFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(\ACK64/$1N2275 ),
    .CLK(CLK),
    .I(\ACK64/IN ),
    .O(\ACK64- ),
    .RST(GND)
  );
  X_ONE   \ACK64/$1I2276/$1I2220  (
    .O(\ACK64/$1I2276/$1N2216 )
  );
  X_BUF   \ACK64/$1I2276/H  (
    .I(\ACK64/$1I2276/$1N2216 ),
    .O(\ACK64/$1N2275 )
  );
  X_ONE   \ACK64/$1I2306/$1I2220  (
    .O(\ACK64/$1I2306/$1N2216 )
  );
  X_BUF   \ACK64/$1I2306/H  (
    .I(\ACK64/$1I2306/$1N2216 ),
    .O(\ACK64/$1N2307 )
  );
  X_MUX2   \ACK64/$1I2310/O  (
    .IA(\ACK64/$1I2310/M01 ),
    .IB(\ACK64/$1I2310/M23 ),
    .O(\ACK64/IN ),
    .SEL(CFG248)
  );
  X_OR2   \ACK64/$1I2310/M01/$1I38  (
    .I0(\ACK64/$1I2310/M01/M1 ),
    .I1(\ACK64/$1I2310/M01/M0 ),
    .O(\ACK64/$1I2310/M01 )
  );
  X_AND3   \ACK64/$1I2310/M01/$1I31  (
    .I0(\NlwInverterSignal_ACK64/$1I2310/M01/$1I31/I0 ),
    .I1(\ACK64/$1N2307 ),
    .I2(ACK64_I),
    .O(\ACK64/$1I2310/M01/M0 )
  );
  X_AND3   \ACK64/$1I2310/M01/$1I30  (
    .I0(\ACK64/D1_9585 ),
    .I1(\ACK64/$1N2307 ),
    .I2(CFG247),
    .O(\ACK64/$1I2310/M01/M1 )
  );
  X_OR2   \ACK64/$1I2310/M23/$1I38  (
    .I0(\ACK64/$1I2310/M23/M1 ),
    .I1(\ACK64/$1I2310/M23/M0 ),
    .O(\ACK64/$1I2310/M23 )
  );
  X_AND3   \ACK64/$1I2310/M23/$1I31  (
    .I0(\NlwInverterSignal_ACK64/$1I2310/M23/$1I31/I0 ),
    .I1(\ACK64/$1N2307 ),
    .I2(\ACK64/D2_9583 ),
    .O(\ACK64/$1I2310/M23/M0 )
  );
  X_AND3   \ACK64/$1I2310/M23/$1I30  (
    .I0(\ACK64/D3_9584 ),
    .I1(\ACK64/$1N2307 ),
    .I2(CFG247),
    .O(\ACK64/$1I2310/M23/M1 )
  );
  X_BUF   \FRAME/$1I2284  (
    .I(FRAME_I),
    .O(\FRAME/D1_9629 )
  );
  X_BUF   \FRAME/$1I2282  (
    .I(\FRAME/D1_9629 ),
    .O(\FRAME/D2_9627 )
  );
  X_BUF   \FRAME/$1I2281  (
    .I(\FRAME/D2_9627 ),
    .O(\FRAME/D3_9628 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \FRAME/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(FRAME_CE),
    .CLK(CLK),
    .I(\NS_FRAME- ),
    .O(FRAME_O),
    .RST(GND)
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \FRAME/IFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(\FRAME/$1N2275 ),
    .CLK(CLK),
    .I(\FRAME/IN ),
    .O(\FRAME- ),
    .RST(GND)
  );
  X_ONE   \FRAME/$1I2276/$1I2220  (
    .O(\FRAME/$1I2276/$1N2216 )
  );
  X_BUF   \FRAME/$1I2276/H  (
    .I(\FRAME/$1I2276/$1N2216 ),
    .O(\FRAME/$1N2275 )
  );
  X_ONE   \FRAME/$1I2306/$1I2220  (
    .O(\FRAME/$1I2306/$1N2216 )
  );
  X_BUF   \FRAME/$1I2306/H  (
    .I(\FRAME/$1I2306/$1N2216 ),
    .O(\FRAME/$1N2307 )
  );
  X_MUX2   \FRAME/$1I2310/O  (
    .IA(\FRAME/$1I2310/M01 ),
    .IB(\FRAME/$1I2310/M23 ),
    .O(\FRAME/IN ),
    .SEL(CFG248)
  );
  X_OR2   \FRAME/$1I2310/M01/$1I38  (
    .I0(\FRAME/$1I2310/M01/M1 ),
    .I1(\FRAME/$1I2310/M01/M0 ),
    .O(\FRAME/$1I2310/M01 )
  );
  X_AND3   \FRAME/$1I2310/M01/$1I31  (
    .I0(\NlwInverterSignal_FRAME/$1I2310/M01/$1I31/I0 ),
    .I1(\FRAME/$1N2307 ),
    .I2(FRAME_I),
    .O(\FRAME/$1I2310/M01/M0 )
  );
  X_AND3   \FRAME/$1I2310/M01/$1I30  (
    .I0(\FRAME/D1_9629 ),
    .I1(\FRAME/$1N2307 ),
    .I2(CFG247),
    .O(\FRAME/$1I2310/M01/M1 )
  );
  X_OR2   \FRAME/$1I2310/M23/$1I38  (
    .I0(\FRAME/$1I2310/M23/M1 ),
    .I1(\FRAME/$1I2310/M23/M0 ),
    .O(\FRAME/$1I2310/M23 )
  );
  X_AND3   \FRAME/$1I2310/M23/$1I31  (
    .I0(\NlwInverterSignal_FRAME/$1I2310/M23/$1I31/I0 ),
    .I1(\FRAME/$1N2307 ),
    .I2(\FRAME/D2_9627 ),
    .O(\FRAME/$1I2310/M23/M0 )
  );
  X_AND3   \FRAME/$1I2310/M23/$1I30  (
    .I0(\FRAME/D3_9628 ),
    .I1(\FRAME/$1N2307 ),
    .I2(CFG247),
    .O(\FRAME/$1I2310/M23/M1 )
  );
  X_ZERO   \$6I1174/$1I2218  (
    .O(\$6I1174/$1N2216 )
  );
  X_BUF   \$6I1174/L  (
    .I(\$6I1174/$1N2216 ),
    .O(\$6N1173 )
  );
  X_BUF   \TRDY/$1I2284  (
    .I(TRDY_I),
    .O(\TRDY/D1_9675 )
  );
  X_BUF   \TRDY/$1I2282  (
    .I(\TRDY/D1_9675 ),
    .O(\TRDY/D2_9673 )
  );
  X_BUF   \TRDY/$1I2281  (
    .I(\TRDY/D2_9673 ),
    .O(\TRDY/D3_9674 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \TRDY/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(TRDY_CE),
    .CLK(CLK),
    .I(\NS_TRDY- ),
    .O(TRDY_O),
    .RST(GND)
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \TRDY/IFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(\TRDY/$1N2275 ),
    .CLK(CLK),
    .I(\TRDY/IN ),
    .O(\TRDY- ),
    .RST(GND)
  );
  X_ONE   \TRDY/$1I2276/$1I2220  (
    .O(\TRDY/$1I2276/$1N2216 )
  );
  X_BUF   \TRDY/$1I2276/H  (
    .I(\TRDY/$1I2276/$1N2216 ),
    .O(\TRDY/$1N2275 )
  );
  X_ONE   \TRDY/$1I2306/$1I2220  (
    .O(\TRDY/$1I2306/$1N2216 )
  );
  X_BUF   \TRDY/$1I2306/H  (
    .I(\TRDY/$1I2306/$1N2216 ),
    .O(\TRDY/$1N2307 )
  );
  X_MUX2   \TRDY/$1I2310/O  (
    .IA(\TRDY/$1I2310/M01 ),
    .IB(\TRDY/$1I2310/M23 ),
    .O(\TRDY/IN ),
    .SEL(CFG248)
  );
  X_OR2   \TRDY/$1I2310/M01/$1I38  (
    .I0(\TRDY/$1I2310/M01/M1 ),
    .I1(\TRDY/$1I2310/M01/M0 ),
    .O(\TRDY/$1I2310/M01 )
  );
  X_AND3   \TRDY/$1I2310/M01/$1I31  (
    .I0(\NlwInverterSignal_TRDY/$1I2310/M01/$1I31/I0 ),
    .I1(\TRDY/$1N2307 ),
    .I2(TRDY_I),
    .O(\TRDY/$1I2310/M01/M0 )
  );
  X_AND3   \TRDY/$1I2310/M01/$1I30  (
    .I0(\TRDY/D1_9675 ),
    .I1(\TRDY/$1N2307 ),
    .I2(CFG247),
    .O(\TRDY/$1I2310/M01/M1 )
  );
  X_OR2   \TRDY/$1I2310/M23/$1I38  (
    .I0(\TRDY/$1I2310/M23/M1 ),
    .I1(\TRDY/$1I2310/M23/M0 ),
    .O(\TRDY/$1I2310/M23 )
  );
  X_AND3   \TRDY/$1I2310/M23/$1I31  (
    .I0(\NlwInverterSignal_TRDY/$1I2310/M23/$1I31/I0 ),
    .I1(\TRDY/$1N2307 ),
    .I2(\TRDY/D2_9673 ),
    .O(\TRDY/$1I2310/M23/M0 )
  );
  X_AND3   \TRDY/$1I2310/M23/$1I30  (
    .I0(\TRDY/D3_9674 ),
    .I1(\TRDY/$1N2307 ),
    .I2(CFG247),
    .O(\TRDY/$1I2310/M23/M1 )
  );
  X_BUF   \REQ64/$1I2284  (
    .I(REQ64_I),
    .O(\REQ64/D1_9719 )
  );
  X_BUF   \REQ64/$1I2282  (
    .I(\REQ64/D1_9719 ),
    .O(\REQ64/D2_9717 )
  );
  X_BUF   \REQ64/$1I2281  (
    .I(\REQ64/D2_9717 ),
    .O(\REQ64/D3_9718 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \REQ64/OFD  (
    .SET(\$6N1173 ),
    .CE(REQ64_CE),
    .CLK(CLK),
    .I(\NS_REQ64- ),
    .O(REQ64_O),
    .RST(GND)
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \REQ64/IFD  (
    .SET(\$6N1173 ),
    .CE(\REQ64/$1N2275 ),
    .CLK(CLK),
    .I(\REQ64/IN ),
    .O(\REQ64- ),
    .RST(GND)
  );
  X_ONE   \REQ64/$1I2276/$1I2220  (
    .O(\REQ64/$1I2276/$1N2216 )
  );
  X_BUF   \REQ64/$1I2276/H  (
    .I(\REQ64/$1I2276/$1N2216 ),
    .O(\REQ64/$1N2275 )
  );
  X_ONE   \REQ64/$1I2306/$1I2220  (
    .O(\REQ64/$1I2306/$1N2216 )
  );
  X_BUF   \REQ64/$1I2306/H  (
    .I(\REQ64/$1I2306/$1N2216 ),
    .O(\REQ64/$1N2307 )
  );
  X_MUX2   \REQ64/$1I2310/O  (
    .IA(\REQ64/$1I2310/M01 ),
    .IB(\REQ64/$1I2310/M23 ),
    .O(\REQ64/IN ),
    .SEL(CFG248)
  );
  X_OR2   \REQ64/$1I2310/M01/$1I38  (
    .I0(\REQ64/$1I2310/M01/M1 ),
    .I1(\REQ64/$1I2310/M01/M0 ),
    .O(\REQ64/$1I2310/M01 )
  );
  X_AND3   \REQ64/$1I2310/M01/$1I31  (
    .I0(\NlwInverterSignal_REQ64/$1I2310/M01/$1I31/I0 ),
    .I1(\REQ64/$1N2307 ),
    .I2(REQ64_I),
    .O(\REQ64/$1I2310/M01/M0 )
  );
  X_AND3   \REQ64/$1I2310/M01/$1I30  (
    .I0(\REQ64/D1_9719 ),
    .I1(\REQ64/$1N2307 ),
    .I2(CFG247),
    .O(\REQ64/$1I2310/M01/M1 )
  );
  X_OR2   \REQ64/$1I2310/M23/$1I38  (
    .I0(\REQ64/$1I2310/M23/M1 ),
    .I1(\REQ64/$1I2310/M23/M0 ),
    .O(\REQ64/$1I2310/M23 )
  );
  X_AND3   \REQ64/$1I2310/M23/$1I31  (
    .I0(\NlwInverterSignal_REQ64/$1I2310/M23/$1I31/I0 ),
    .I1(\REQ64/$1N2307 ),
    .I2(\REQ64/D2_9717 ),
    .O(\REQ64/$1I2310/M23/M0 )
  );
  X_AND3   \REQ64/$1I2310/M23/$1I30  (
    .I0(\REQ64/D3_9718 ),
    .I1(\REQ64/$1N2307 ),
    .I2(CFG247),
    .O(\REQ64/$1I2310/M23/M1 )
  );
  X_BUF   \IRDY/$1I2284  (
    .I(IRDY_I),
    .O(\IRDY/D1_9763 )
  );
  X_BUF   \IRDY/$1I2282  (
    .I(\IRDY/D1_9763 ),
    .O(\IRDY/D2_9761 )
  );
  X_BUF   \IRDY/$1I2281  (
    .I(\IRDY/D2_9761 ),
    .O(\IRDY/D3_9762 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \IRDY/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(IRDY_CE),
    .CLK(CLK),
    .I(\NS_IRDY- ),
    .O(IRDY_O),
    .RST(GND)
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \IRDY/IFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(\IRDY/$1N2275 ),
    .CLK(CLK),
    .I(\IRDY/IN ),
    .O(\IRDY- ),
    .RST(GND)
  );
  X_ONE   \IRDY/$1I2276/$1I2220  (
    .O(\IRDY/$1I2276/$1N2216 )
  );
  X_BUF   \IRDY/$1I2276/H  (
    .I(\IRDY/$1I2276/$1N2216 ),
    .O(\IRDY/$1N2275 )
  );
  X_ONE   \IRDY/$1I2306/$1I2220  (
    .O(\IRDY/$1I2306/$1N2216 )
  );
  X_BUF   \IRDY/$1I2306/H  (
    .I(\IRDY/$1I2306/$1N2216 ),
    .O(\IRDY/$1N2307 )
  );
  X_MUX2   \IRDY/$1I2310/O  (
    .IA(\IRDY/$1I2310/M01 ),
    .IB(\IRDY/$1I2310/M23 ),
    .O(\IRDY/IN ),
    .SEL(CFG248)
  );
  X_OR2   \IRDY/$1I2310/M01/$1I38  (
    .I0(\IRDY/$1I2310/M01/M1 ),
    .I1(\IRDY/$1I2310/M01/M0 ),
    .O(\IRDY/$1I2310/M01 )
  );
  X_AND3   \IRDY/$1I2310/M01/$1I31  (
    .I0(\NlwInverterSignal_IRDY/$1I2310/M01/$1I31/I0 ),
    .I1(\IRDY/$1N2307 ),
    .I2(IRDY_I),
    .O(\IRDY/$1I2310/M01/M0 )
  );
  X_AND3   \IRDY/$1I2310/M01/$1I30  (
    .I0(\IRDY/D1_9763 ),
    .I1(\IRDY/$1N2307 ),
    .I2(CFG247),
    .O(\IRDY/$1I2310/M01/M1 )
  );
  X_OR2   \IRDY/$1I2310/M23/$1I38  (
    .I0(\IRDY/$1I2310/M23/M1 ),
    .I1(\IRDY/$1I2310/M23/M0 ),
    .O(\IRDY/$1I2310/M23 )
  );
  X_AND3   \IRDY/$1I2310/M23/$1I31  (
    .I0(\NlwInverterSignal_IRDY/$1I2310/M23/$1I31/I0 ),
    .I1(\IRDY/$1N2307 ),
    .I2(\IRDY/D2_9761 ),
    .O(\IRDY/$1I2310/M23/M0 )
  );
  X_AND3   \IRDY/$1I2310/M23/$1I30  (
    .I0(\IRDY/D3_9762 ),
    .I1(\IRDY/$1N2307 ),
    .I2(CFG247),
    .O(\IRDY/$1I2310/M23/M1 )
  );
  X_BUF   \STOP/$1I2284  (
    .I(STOP_I),
    .O(\STOP/D1_9807 )
  );
  X_BUF   \STOP/$1I2282  (
    .I(\STOP/D1_9807 ),
    .O(\STOP/D2_9805 )
  );
  X_BUF   \STOP/$1I2281  (
    .I(\STOP/D2_9805 ),
    .O(\STOP/D3_9806 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \STOP/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(STOP_CE),
    .CLK(CLK),
    .I(\NS_STOP- ),
    .O(STOP_O),
    .RST(GND)
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \STOP/IFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(\STOP/$1N2275 ),
    .CLK(CLK),
    .I(\STOP/IN ),
    .O(\STOP- ),
    .RST(GND)
  );
  X_ONE   \STOP/$1I2276/$1I2220  (
    .O(\STOP/$1I2276/$1N2216 )
  );
  X_BUF   \STOP/$1I2276/H  (
    .I(\STOP/$1I2276/$1N2216 ),
    .O(\STOP/$1N2275 )
  );
  X_ONE   \STOP/$1I2306/$1I2220  (
    .O(\STOP/$1I2306/$1N2216 )
  );
  X_BUF   \STOP/$1I2306/H  (
    .I(\STOP/$1I2306/$1N2216 ),
    .O(\STOP/$1N2307 )
  );
  X_MUX2   \STOP/$1I2310/O  (
    .IA(\STOP/$1I2310/M01 ),
    .IB(\STOP/$1I2310/M23 ),
    .O(\STOP/IN ),
    .SEL(CFG248)
  );
  X_OR2   \STOP/$1I2310/M01/$1I38  (
    .I0(\STOP/$1I2310/M01/M1 ),
    .I1(\STOP/$1I2310/M01/M0 ),
    .O(\STOP/$1I2310/M01 )
  );
  X_AND3   \STOP/$1I2310/M01/$1I31  (
    .I0(\NlwInverterSignal_STOP/$1I2310/M01/$1I31/I0 ),
    .I1(\STOP/$1N2307 ),
    .I2(STOP_I),
    .O(\STOP/$1I2310/M01/M0 )
  );
  X_AND3   \STOP/$1I2310/M01/$1I30  (
    .I0(\STOP/D1_9807 ),
    .I1(\STOP/$1N2307 ),
    .I2(CFG247),
    .O(\STOP/$1I2310/M01/M1 )
  );
  X_OR2   \STOP/$1I2310/M23/$1I38  (
    .I0(\STOP/$1I2310/M23/M1 ),
    .I1(\STOP/$1I2310/M23/M0 ),
    .O(\STOP/$1I2310/M23 )
  );
  X_AND3   \STOP/$1I2310/M23/$1I31  (
    .I0(\NlwInverterSignal_STOP/$1I2310/M23/$1I31/I0 ),
    .I1(\STOP/$1N2307 ),
    .I2(\STOP/D2_9805 ),
    .O(\STOP/$1I2310/M23/M0 )
  );
  X_AND3   \STOP/$1I2310/M23/$1I30  (
    .I0(\STOP/D3_9806 ),
    .I1(\STOP/$1N2307 ),
    .I2(CFG247),
    .O(\STOP/$1I2310/M23/M1 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PERR/IFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(\PERR/$1N2286 ),
    .CLK(CLK),
    .I(PERR_I),
    .O(\PERR- ),
    .RST(GND)
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PERR/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(\PERR/$1N2289 ),
    .CLK(CLK),
    .I(\NS_PERR- ),
    .O(PERR_O),
    .RST(GND)
  );
  X_ONE   \PERR/$1I2285/$1I2220  (
    .O(\PERR/$1I2285/$1N2216 )
  );
  X_BUF   \PERR/$1I2285/H  (
    .I(\PERR/$1I2285/$1N2216 ),
    .O(\PERR/$1N2286 )
  );
  X_ONE   \PERR/$1I2288/$1I2220  (
    .O(\PERR/$1I2288/$1N2216 )
  );
  X_BUF   \PERR/$1I2288/H  (
    .I(\PERR/$1I2288/$1N2216 ),
    .O(\PERR/$1N2289 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \SERR/IFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(\SERR/$1N2286 ),
    .CLK(CLK),
    .I(SERR_I),
    .O(\SERR- ),
    .RST(GND)
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \SERR/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(\SERR/$1N2289 ),
    .CLK(CLK),
    .I(\NS_SERR- ),
    .O(SERR_O),
    .RST(GND)
  );
  X_ONE   \SERR/$1I2285/$1I2220  (
    .O(\SERR/$1I2285/$1N2216 )
  );
  X_BUF   \SERR/$1I2285/H  (
    .I(\SERR/$1I2285/$1N2216 ),
    .O(\SERR/$1N2286 )
  );
  X_ONE   \SERR/$1I2288/$1I2220  (
    .O(\SERR/$1I2288/$1N2216 )
  );
  X_BUF   \SERR/$1I2288/H  (
    .I(\SERR/$1I2288/$1N2216 ),
    .O(\SERR/$1N2289 )
  );
  X_ZERO   \$6I950/$1I2218  (
    .O(\$6I950/$1N2216 )
  );
  X_BUF   \$6I950/L  (
    .I(\$6I950/$1N2216 ),
    .O(\NS_SERR- )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \IDSEL/IFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(\IDSEL/$1N2286 ),
    .CLK(CLK),
    .I(IDSEL_IN),
    .O(IDSEL),
    .RST(GND)
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \IDSEL/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(\IDSEL/$1N2289 ),
    .CLK(CLK),
    .I(NS_IDSEL),
    .O(IDSEL_O),
    .RST(GND)
  );
  X_ONE   \IDSEL/$1I2285/$1I2220  (
    .O(\IDSEL/$1I2285/$1N2216 )
  );
  X_BUF   \IDSEL/$1I2285/H  (
    .I(\IDSEL/$1I2285/$1N2216 ),
    .O(\IDSEL/$1N2286 )
  );
  X_ONE   \IDSEL/$1I2288/$1I2220  (
    .O(\IDSEL/$1I2288/$1N2216 )
  );
  X_BUF   \IDSEL/$1I2288/H  (
    .I(\IDSEL/$1I2288/$1N2216 ),
    .O(\IDSEL/$1N2289 )
  );
  X_ZERO   \$6I961/$1I2218  (
    .O(\$6I961/$1N2216 )
  );
  X_BUF   \$6I961/L  (
    .I(\$6I961/$1N2216 ),
    .O(NS_IDSEL)
  );
  X_AND2   \$7I576/$1I9  (
    .I0(INTACK),
    .I1(CFG240),
    .O(\$7I576/M1 )
  );
  X_OR2   \$7I576/$1I8  (
    .I0(\$7I576/M1 ),
    .I1(\$7I576/M0 ),
    .O(NS_BASE_HIT2)
  );
  X_AND2   \$7I576/$1I7  (
    .I0(\NlwInverterSignal_$7I576/$1I7/I0 ),
    .I1(NS_BASE_HIT2_INT),
    .O(\$7I576/M0 )
  );
  X_AND2   \$7I577/$1I9  (
    .I0(INTACKQ),
    .I1(CFG240),
    .O(\$7I577/M1 )
  );
  X_OR2   \$7I577/$1I8  (
    .I0(\$7I577/M1 ),
    .I1(\$7I577/M0 ),
    .O(NlwRenamedSig_OI_BASE_HIT2)
  );
  X_AND2   \$7I577/$1I7  (
    .I0(\NlwInverterSignal_$7I577/$1I7/I0 ),
    .I1(BASE_HIT2_INT),
    .O(\$7I577/M0 )
  );
  X_AND4   \$7I580/AND4  (
    .I0(\$7I580/$1N2275 ),
    .I1(\$7I580/$1N2276 ),
    .I2(\$7I580/$1N2277 ),
    .I3(\$7I580/$1N2283 ),
    .O(\$7N583 )
  );
  X_INV   \$7I580/INV3  (
    .I(NlwRenamedSig_OI_S_CBE3),
    .O(\$7I580/$1N2283 )
  );
  X_INV   \$7I580/INV2  (
    .I(NlwRenamedSig_OI_S_CBE2),
    .O(\$7I580/$1N2277 )
  );
  X_INV   \$7I580/INV1  (
    .I(NlwRenamedSig_OI_S_CBE1),
    .O(\$7I580/$1N2276 )
  );
  X_INV   \$7I580/INV0  (
    .I(NlwRenamedSig_OI_S_CBE0),
    .O(\$7I580/$1N2275 )
  );
  X_AND2   \$7I622/$1I9  (
    .I0(\$7N625 ),
    .I1(CFG240),
    .O(\$7I622/M1 )
  );
  X_OR2   \$7I622/$1I8  (
    .I0(\$7I622/M1 ),
    .I1(\$7I622/M0 ),
    .O(NS_BH64_2)
  );
  X_AND2   \$7I622/$1I7  (
    .I0(\NlwInverterSignal_$7I622/$1I7/I0 ),
    .I1(NS_BH64_2_INT),
    .O(\$7I622/M0 )
  );
  X_AND2   \$7I623/$1I9  (
    .I0(\$7N621 ),
    .I1(CFG240),
    .O(\$7I623/M1 )
  );
  X_OR2   \$7I623/$1I8  (
    .I0(\$7I623/M1 ),
    .I1(\$7I623/M0 ),
    .O(BH64_2)
  );
  X_AND2   \$7I623/$1I7  (
    .I0(\NlwInverterSignal_$7I623/$1I7/I0 ),
    .I1(BH64_2_INT),
    .O(\$7I623/M0 )
  );
  X_ZERO   \$7I632/$1I2218  (
    .O(\$7I632/$1N2216 )
  );
  X_BUF   \$7I632/L  (
    .I(\$7I632/$1N2216 ),
    .O(\$7N625 )
  );
  X_ZERO   \$7I633/$1I2218  (
    .O(\$7I633/$1N2216 )
  );
  X_BUF   \$7I633/L  (
    .I(\$7I633/$1N2216 ),
    .O(\$7N621 )
  );
  X_ZERO   \$7I746/$1I2218  (
    .O(\$7I746/$1N2216 )
  );
  X_BUF   \$7I746/L  (
    .I(\$7I746/$1N2216 ),
    .O(\$7N745 )
  );
  X_AND2   \$7I824/$1I9  (
    .I0(NlwRenamedSig_OI_OE_ADO_LB),
    .I1(CFG255),
    .O(\$7I824/M1 )
  );
  X_OR2   \$7I824/$1I8  (
    .I0(\$7I824/M1 ),
    .I1(\$7I824/M0 ),
    .O(NlwRenamedSig_OI_CSR32)
  );
  X_AND2   \$7I824/$1I7  (
    .I0(\NlwInverterSignal_$7I824/$1I7/I0 ),
    .I1(\$7N147 ),
    .O(\$7I824/M0 )
  );
  X_AND2   \$7I826/$1I9  (
    .I0(NlwRenamedSig_OI_OE_CBE),
    .I1(CFG255),
    .O(\$7I826/M1 )
  );
  X_OR2   \$7I826/$1I8  (
    .I0(\$7I826/M1 ),
    .I1(\$7I826/M0 ),
    .O(NlwRenamedSig_OI_CSR33)
  );
  X_AND2   \$7I826/$1I7  (
    .I0(\NlwInverterSignal_$7I826/$1I7/I0 ),
    .I1(\$7N148 ),
    .O(\$7I826/M0 )
  );
  X_AND2   \$7I828/$1I9  (
    .I0(NlwRenamedSig_OI_OE_PAR),
    .I1(CFG255),
    .O(\$7I828/M1 )
  );
  X_OR2   \$7I828/$1I8  (
    .I0(\$7I828/M1 ),
    .I1(\$7I828/M0 ),
    .O(NlwRenamedSig_OI_CSR34)
  );
  X_AND2   \$7I828/$1I7  (
    .I0(\NlwInverterSignal_$7I828/$1I7/I0 ),
    .I1(\$7N149 ),
    .O(\$7I828/M0 )
  );
  X_AND2   \$7I830/$1I9  (
    .I0(\$7N855 ),
    .I1(CFG255),
    .O(\$7I830/M1 )
  );
  X_OR2   \$7I830/$1I8  (
    .I0(\$7I830/M1 ),
    .I1(\$7I830/M0 ),
    .O(NlwRenamedSig_OI_CSR35)
  );
  X_AND2   \$7I830/$1I7  (
    .I0(\NlwInverterSignal_$7I830/$1I7/I0 ),
    .I1(\$7N152 ),
    .O(\$7I830/M0 )
  );
  X_AND2   \$7I832/$1I9  (
    .I0(NlwRenamedSig_OI_OE_ADO_LB64),
    .I1(CFG255),
    .O(\$7I832/M1 )
  );
  X_OR2   \$7I832/$1I8  (
    .I0(\$7I832/M1 ),
    .I1(\$7I832/M0 ),
    .O(NlwRenamedSig_OI_CSR36)
  );
  X_AND2   \$7I832/$1I7  (
    .I0(\NlwInverterSignal_$7I832/$1I7/I0 ),
    .I1(\$7N156 ),
    .O(\$7I832/M0 )
  );
  X_AND2   \$7I834/$1I9  (
    .I0(NlwRenamedSig_OI_OE_CBE64),
    .I1(CFG255),
    .O(\$7I834/M1 )
  );
  X_OR2   \$7I834/$1I8  (
    .I0(\$7I834/M1 ),
    .I1(\$7I834/M0 ),
    .O(NlwRenamedSig_OI_CSR37)
  );
  X_AND2   \$7I834/$1I7  (
    .I0(\NlwInverterSignal_$7I834/$1I7/I0 ),
    .I1(\$7N160 ),
    .O(\$7I834/M0 )
  );
  X_AND2   \$7I836/$1I9  (
    .I0(NlwRenamedSig_OI_OE_PAR64),
    .I1(CFG255),
    .O(\$7I836/M1 )
  );
  X_OR2   \$7I836/$1I8  (
    .I0(\$7I836/M1 ),
    .I1(\$7I836/M0 ),
    .O(NlwRenamedSig_OI_CSR38)
  );
  X_AND2   \$7I836/$1I7  (
    .I0(\NlwInverterSignal_$7I836/$1I7/I0 ),
    .I1(\$7N163 ),
    .O(\$7I836/M0 )
  );
  X_AND2   \$7I838/$1I9  (
    .I0(\$7N859 ),
    .I1(CFG255),
    .O(\$7I838/M1 )
  );
  X_OR2   \$7I838/$1I8  (
    .I0(\$7I838/M1 ),
    .I1(\$7I838/M0 ),
    .O(NlwRenamedSig_OI_CSR39)
  );
  X_AND2   \$7I838/$1I7  (
    .I0(\NlwInverterSignal_$7I838/$1I7/I0 ),
    .I1(SET13),
    .O(\$7I838/M0 )
  );
  X_ONE   \$7I861/$1I2220  (
    .O(\$7I861/$1N2216 )
  );
  X_BUF   \$7I861/H  (
    .I(\$7I861/$1N2216 ),
    .O(\$7N855 )
  );
  X_ONE   \$7I862/$1I2220  (
    .O(\$7I862/$1N2216 )
  );
  X_BUF   \$7I862/H  (
    .I(\$7I862/$1N2216 ),
    .O(\$7N859 )
  );
  X_AND2   \PCI-CBE/$1I2773  (
    .I0(\NlwInverterSignal_PCI-CBE/$1I2773/I0 ),
    .I1(ATTEMPT64),
    .O(\PCI-CBE/SWITCH )
  );
  X_AND2   \PCI-CBE/IO3/$1I2316  (
    .I0(\PCI-CBE/TO_ACK ),
    .I1(\PCI-CBE/TO_SW ),
    .O(\PCI-CBE/IO3/$1N2321 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-CBE/IO3/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(CBEOUT3),
    .O(CBE_O3),
    .RST(GND)
  );
  X_AND2   \PCI-CBE/IO3/$1I2296/$1I9  (
    .I0(SHADOW_CBE3),
    .I1(OUT_SEL),
    .O(\PCI-CBE/IO3/$1I2296/M1 )
  );
  X_OR2   \PCI-CBE/IO3/$1I2296/$1I8  (
    .I0(\PCI-CBE/IO3/$1I2296/M1 ),
    .I1(\PCI-CBE/IO3/$1I2296/M0 ),
    .O(\PCI-CBE/IO3/D_SLO )
  );
  X_AND2   \PCI-CBE/IO3/$1I2296/$1I7  (
    .I0(\NlwInverterSignal_PCI-CBE/IO3/$1I2296/$1I7/I0 ),
    .I1(M_CBE_INT3),
    .O(\PCI-CBE/IO3/$1I2296/M0 )
  );
  X_AND2   \PCI-CBE/IO3/$1I2303/$1I9  (
    .I0(FAIL_CBH7),
    .I1(\PCI-CBE/IO3/$1N2321 ),
    .O(\PCI-CBE/IO3/$1I2303/M1 )
  );
  X_OR2   \PCI-CBE/IO3/$1I2303/$1I8  (
    .I0(\PCI-CBE/IO3/$1I2303/M1 ),
    .I1(\PCI-CBE/IO3/$1I2303/M0 ),
    .O(CBEOUT3)
  );
  X_AND2   \PCI-CBE/IO3/$1I2303/$1I7  (
    .I0(\NlwInverterSignal_PCI-CBE/IO3/$1I2303/$1I7/I0 ),
    .I1(\PCI-CBE/IO3/D_SLO ),
    .O(\PCI-CBE/IO3/$1I2303/M0 )
  );
  X_AND2   \PCI-CBE/IO2/$1I2316  (
    .I0(\PCI-CBE/TO_ACK ),
    .I1(\PCI-CBE/TO_SW ),
    .O(\PCI-CBE/IO2/$1N2321 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-CBE/IO2/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(CBEOUT2),
    .O(CBE_O2),
    .RST(GND)
  );
  X_AND2   \PCI-CBE/IO2/$1I2296/$1I9  (
    .I0(SHADOW_CBE2),
    .I1(OUT_SEL),
    .O(\PCI-CBE/IO2/$1I2296/M1 )
  );
  X_OR2   \PCI-CBE/IO2/$1I2296/$1I8  (
    .I0(\PCI-CBE/IO2/$1I2296/M1 ),
    .I1(\PCI-CBE/IO2/$1I2296/M0 ),
    .O(\PCI-CBE/IO2/D_SLO )
  );
  X_AND2   \PCI-CBE/IO2/$1I2296/$1I7  (
    .I0(\NlwInverterSignal_PCI-CBE/IO2/$1I2296/$1I7/I0 ),
    .I1(M_CBE_INT2),
    .O(\PCI-CBE/IO2/$1I2296/M0 )
  );
  X_AND2   \PCI-CBE/IO2/$1I2303/$1I9  (
    .I0(FAIL_CBH6),
    .I1(\PCI-CBE/IO2/$1N2321 ),
    .O(\PCI-CBE/IO2/$1I2303/M1 )
  );
  X_OR2   \PCI-CBE/IO2/$1I2303/$1I8  (
    .I0(\PCI-CBE/IO2/$1I2303/M1 ),
    .I1(\PCI-CBE/IO2/$1I2303/M0 ),
    .O(CBEOUT2)
  );
  X_AND2   \PCI-CBE/IO2/$1I2303/$1I7  (
    .I0(\NlwInverterSignal_PCI-CBE/IO2/$1I2303/$1I7/I0 ),
    .I1(\PCI-CBE/IO2/D_SLO ),
    .O(\PCI-CBE/IO2/$1I2303/M0 )
  );
  X_AND2   \PCI-CBE/IO1/$1I2316  (
    .I0(\PCI-CBE/TO_ACK ),
    .I1(\PCI-CBE/TO_SW ),
    .O(\PCI-CBE/IO1/$1N2321 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-CBE/IO1/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(CBEOUT1),
    .O(CBE_O1),
    .RST(GND)
  );
  X_AND2   \PCI-CBE/IO1/$1I2296/$1I9  (
    .I0(SHADOW_CBE1),
    .I1(OUT_SEL),
    .O(\PCI-CBE/IO1/$1I2296/M1 )
  );
  X_OR2   \PCI-CBE/IO1/$1I2296/$1I8  (
    .I0(\PCI-CBE/IO1/$1I2296/M1 ),
    .I1(\PCI-CBE/IO1/$1I2296/M0 ),
    .O(\PCI-CBE/IO1/D_SLO )
  );
  X_AND2   \PCI-CBE/IO1/$1I2296/$1I7  (
    .I0(\NlwInverterSignal_PCI-CBE/IO1/$1I2296/$1I7/I0 ),
    .I1(M_CBE_INT1),
    .O(\PCI-CBE/IO1/$1I2296/M0 )
  );
  X_AND2   \PCI-CBE/IO1/$1I2303/$1I9  (
    .I0(FAIL_CBH5),
    .I1(\PCI-CBE/IO1/$1N2321 ),
    .O(\PCI-CBE/IO1/$1I2303/M1 )
  );
  X_OR2   \PCI-CBE/IO1/$1I2303/$1I8  (
    .I0(\PCI-CBE/IO1/$1I2303/M1 ),
    .I1(\PCI-CBE/IO1/$1I2303/M0 ),
    .O(CBEOUT1)
  );
  X_AND2   \PCI-CBE/IO1/$1I2303/$1I7  (
    .I0(\NlwInverterSignal_PCI-CBE/IO1/$1I2303/$1I7/I0 ),
    .I1(\PCI-CBE/IO1/D_SLO ),
    .O(\PCI-CBE/IO1/$1I2303/M0 )
  );
  X_AND2   \PCI-CBE/IO0/$1I2316  (
    .I0(\PCI-CBE/TO_ACK ),
    .I1(\PCI-CBE/TO_SW ),
    .O(\PCI-CBE/IO0/$1N2321 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-CBE/IO0/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(CBEOUT0),
    .O(CBE_O0),
    .RST(GND)
  );
  X_AND2   \PCI-CBE/IO0/$1I2296/$1I9  (
    .I0(SHADOW_CBE0),
    .I1(OUT_SEL),
    .O(\PCI-CBE/IO0/$1I2296/M1 )
  );
  X_OR2   \PCI-CBE/IO0/$1I2296/$1I8  (
    .I0(\PCI-CBE/IO0/$1I2296/M1 ),
    .I1(\PCI-CBE/IO0/$1I2296/M0 ),
    .O(\PCI-CBE/IO0/D_SLO )
  );
  X_AND2   \PCI-CBE/IO0/$1I2296/$1I7  (
    .I0(\NlwInverterSignal_PCI-CBE/IO0/$1I2296/$1I7/I0 ),
    .I1(M_CBE_INT0),
    .O(\PCI-CBE/IO0/$1I2296/M0 )
  );
  X_AND2   \PCI-CBE/IO0/$1I2303/$1I9  (
    .I0(FAIL_CBH4),
    .I1(\PCI-CBE/IO0/$1N2321 ),
    .O(\PCI-CBE/IO0/$1I2303/M1 )
  );
  X_OR2   \PCI-CBE/IO0/$1I2303/$1I8  (
    .I0(\PCI-CBE/IO0/$1I2303/M1 ),
    .I1(\PCI-CBE/IO0/$1I2303/M0 ),
    .O(CBEOUT0)
  );
  X_AND2   \PCI-CBE/IO0/$1I2303/$1I7  (
    .I0(\NlwInverterSignal_PCI-CBE/IO0/$1I2303/$1I7/I0 ),
    .I1(\PCI-CBE/IO0/D_SLO ),
    .O(\PCI-CBE/IO0/$1I2303/M0 )
  );
  X_AND2   \PCI-CBE/$1I2777/$1I9  (
    .I0(\PCI-CBE/SWITCH ),
    .I1(CFG253),
    .O(\PCI-CBE/$1I2777/M1 )
  );
  X_OR2   \PCI-CBE/$1I2777/$1I8  (
    .I0(\PCI-CBE/$1I2777/M1 ),
    .I1(\PCI-CBE/$1I2777/M0 ),
    .O(\PCI-CBE/TO_SW )
  );
  X_AND2   \PCI-CBE/$1I2777/$1I7  (
    .I0(\NlwInverterSignal_PCI-CBE/$1I2777/$1I7/I0 ),
    .I1(FAIL64_INT),
    .O(\PCI-CBE/$1I2777/M0 )
  );
  X_AND2   \PCI-CBE/$1I2779/$1I9  (
    .I0(ACK64_I),
    .I1(CFG253),
    .O(\PCI-CBE/$1I2779/M1 )
  );
  X_OR2   \PCI-CBE/$1I2779/$1I8  (
    .I0(\PCI-CBE/$1I2779/M1 ),
    .I1(\PCI-CBE/$1I2779/M0 ),
    .O(\PCI-CBE/TO_ACK )
  );
  X_AND2   \PCI-CBE/$1I2779/$1I7  (
    .I0(\NlwInverterSignal_PCI-CBE/$1I2779/$1I7/I0 ),
    .I1(\PCI-CBE/$1N2786 ),
    .O(\PCI-CBE/$1I2779/M0 )
  );
  X_ONE   \PCI-CBE/$1I2787/$1I2220  (
    .O(\PCI-CBE/$1I2787/$1N2216 )
  );
  X_BUF   \PCI-CBE/$1I2787/H  (
    .I(\PCI-CBE/$1I2787/$1N2216 ),
    .O(\PCI-CBE/$1N2786 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD/IO28/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT28),
    .O(AD_O28),
    .RST(GND)
  );
  X_AND2   \PCI-AD/IO28/$1I2246/$1I9  (
    .I0(FAIL_ADH60),
    .I1(FAIL64_INT),
    .O(\PCI-AD/IO28/$1I2246/M1 )
  );
  X_OR2   \PCI-AD/IO28/$1I2246/$1I8  (
    .I0(\PCI-AD/IO28/$1I2246/M1 ),
    .I1(\PCI-AD/IO28/$1I2246/M0 ),
    .O(ADOUT28)
  );
  X_AND2   \PCI-AD/IO28/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/IO28/$1I2246/$1I7/I0 ),
    .I1(\PCI-AD/D_SLO28 ),
    .O(\PCI-AD/IO28/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD/IO30/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT30),
    .O(AD_O30),
    .RST(GND)
  );
  X_AND2   \PCI-AD/IO30/$1I2246/$1I9  (
    .I0(FAIL_ADH62),
    .I1(FAIL64_INT),
    .O(\PCI-AD/IO30/$1I2246/M1 )
  );
  X_OR2   \PCI-AD/IO30/$1I2246/$1I8  (
    .I0(\PCI-AD/IO30/$1I2246/M1 ),
    .I1(\PCI-AD/IO30/$1I2246/M0 ),
    .O(ADOUT30)
  );
  X_AND2   \PCI-AD/IO30/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/IO30/$1I2246/$1I7/I0 ),
    .I1(\PCI-AD/D_SLO30 ),
    .O(\PCI-AD/IO30/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD/IO29/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT29),
    .O(AD_O29),
    .RST(GND)
  );
  X_AND2   \PCI-AD/IO29/$1I2246/$1I9  (
    .I0(FAIL_ADH61),
    .I1(FAIL64_INT),
    .O(\PCI-AD/IO29/$1I2246/M1 )
  );
  X_OR2   \PCI-AD/IO29/$1I2246/$1I8  (
    .I0(\PCI-AD/IO29/$1I2246/M1 ),
    .I1(\PCI-AD/IO29/$1I2246/M0 ),
    .O(ADOUT29)
  );
  X_AND2   \PCI-AD/IO29/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/IO29/$1I2246/$1I7/I0 ),
    .I1(\PCI-AD/D_SLO29 ),
    .O(\PCI-AD/IO29/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD/IO31/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT31),
    .O(AD_O31),
    .RST(GND)
  );
  X_AND2   \PCI-AD/IO31/$1I2246/$1I9  (
    .I0(FAIL_ADH63),
    .I1(FAIL64_INT),
    .O(\PCI-AD/IO31/$1I2246/M1 )
  );
  X_OR2   \PCI-AD/IO31/$1I2246/$1I8  (
    .I0(\PCI-AD/IO31/$1I2246/M1 ),
    .I1(\PCI-AD/IO31/$1I2246/M0 ),
    .O(ADOUT31)
  );
  X_AND2   \PCI-AD/IO31/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/IO31/$1I2246/$1I7/I0 ),
    .I1(\PCI-AD/D_SLO31 ),
    .O(\PCI-AD/IO31/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD/IO20/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT20),
    .O(AD_O20),
    .RST(GND)
  );
  X_AND2   \PCI-AD/IO20/$1I2246/$1I9  (
    .I0(FAIL_ADH52),
    .I1(FAIL64_INT),
    .O(\PCI-AD/IO20/$1I2246/M1 )
  );
  X_OR2   \PCI-AD/IO20/$1I2246/$1I8  (
    .I0(\PCI-AD/IO20/$1I2246/M1 ),
    .I1(\PCI-AD/IO20/$1I2246/M0 ),
    .O(ADOUT20)
  );
  X_AND2   \PCI-AD/IO20/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/IO20/$1I2246/$1I7/I0 ),
    .I1(\PCI-AD/D_SLO20 ),
    .O(\PCI-AD/IO20/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD/IO22/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT22),
    .O(AD_O22),
    .RST(GND)
  );
  X_AND2   \PCI-AD/IO22/$1I2246/$1I9  (
    .I0(FAIL_ADH54),
    .I1(FAIL64_INT),
    .O(\PCI-AD/IO22/$1I2246/M1 )
  );
  X_OR2   \PCI-AD/IO22/$1I2246/$1I8  (
    .I0(\PCI-AD/IO22/$1I2246/M1 ),
    .I1(\PCI-AD/IO22/$1I2246/M0 ),
    .O(ADOUT22)
  );
  X_AND2   \PCI-AD/IO22/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/IO22/$1I2246/$1I7/I0 ),
    .I1(\PCI-AD/D_SLO22 ),
    .O(\PCI-AD/IO22/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD/IO21/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT21),
    .O(AD_O21),
    .RST(GND)
  );
  X_AND2   \PCI-AD/IO21/$1I2246/$1I9  (
    .I0(FAIL_ADH53),
    .I1(FAIL64_INT),
    .O(\PCI-AD/IO21/$1I2246/M1 )
  );
  X_OR2   \PCI-AD/IO21/$1I2246/$1I8  (
    .I0(\PCI-AD/IO21/$1I2246/M1 ),
    .I1(\PCI-AD/IO21/$1I2246/M0 ),
    .O(ADOUT21)
  );
  X_AND2   \PCI-AD/IO21/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/IO21/$1I2246/$1I7/I0 ),
    .I1(\PCI-AD/D_SLO21 ),
    .O(\PCI-AD/IO21/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD/IO23/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT23),
    .O(AD_O23),
    .RST(GND)
  );
  X_AND2   \PCI-AD/IO23/$1I2246/$1I9  (
    .I0(FAIL_ADH55),
    .I1(FAIL64_INT),
    .O(\PCI-AD/IO23/$1I2246/M1 )
  );
  X_OR2   \PCI-AD/IO23/$1I2246/$1I8  (
    .I0(\PCI-AD/IO23/$1I2246/M1 ),
    .I1(\PCI-AD/IO23/$1I2246/M0 ),
    .O(ADOUT23)
  );
  X_AND2   \PCI-AD/IO23/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/IO23/$1I2246/$1I7/I0 ),
    .I1(\PCI-AD/D_SLO23 ),
    .O(\PCI-AD/IO23/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD/IO12/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT12),
    .O(AD_O12),
    .RST(GND)
  );
  X_AND2   \PCI-AD/IO12/$1I2246/$1I9  (
    .I0(FAIL_ADH44),
    .I1(FAIL64_INT),
    .O(\PCI-AD/IO12/$1I2246/M1 )
  );
  X_OR2   \PCI-AD/IO12/$1I2246/$1I8  (
    .I0(\PCI-AD/IO12/$1I2246/M1 ),
    .I1(\PCI-AD/IO12/$1I2246/M0 ),
    .O(ADOUT12)
  );
  X_AND2   \PCI-AD/IO12/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/IO12/$1I2246/$1I7/I0 ),
    .I1(\PCI-AD/D_SLO12 ),
    .O(\PCI-AD/IO12/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD/IO14/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT14),
    .O(AD_O14),
    .RST(GND)
  );
  X_AND2   \PCI-AD/IO14/$1I2246/$1I9  (
    .I0(FAIL_ADH46),
    .I1(FAIL64_INT),
    .O(\PCI-AD/IO14/$1I2246/M1 )
  );
  X_OR2   \PCI-AD/IO14/$1I2246/$1I8  (
    .I0(\PCI-AD/IO14/$1I2246/M1 ),
    .I1(\PCI-AD/IO14/$1I2246/M0 ),
    .O(ADOUT14)
  );
  X_AND2   \PCI-AD/IO14/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/IO14/$1I2246/$1I7/I0 ),
    .I1(\PCI-AD/D_SLO14 ),
    .O(\PCI-AD/IO14/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD/IO13/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT13),
    .O(AD_O13),
    .RST(GND)
  );
  X_AND2   \PCI-AD/IO13/$1I2246/$1I9  (
    .I0(FAIL_ADH45),
    .I1(FAIL64_INT),
    .O(\PCI-AD/IO13/$1I2246/M1 )
  );
  X_OR2   \PCI-AD/IO13/$1I2246/$1I8  (
    .I0(\PCI-AD/IO13/$1I2246/M1 ),
    .I1(\PCI-AD/IO13/$1I2246/M0 ),
    .O(ADOUT13)
  );
  X_AND2   \PCI-AD/IO13/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/IO13/$1I2246/$1I7/I0 ),
    .I1(\PCI-AD/D_SLO13 ),
    .O(\PCI-AD/IO13/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD/IO15/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT15),
    .O(AD_O15),
    .RST(GND)
  );
  X_AND2   \PCI-AD/IO15/$1I2246/$1I9  (
    .I0(FAIL_ADH47),
    .I1(FAIL64_INT),
    .O(\PCI-AD/IO15/$1I2246/M1 )
  );
  X_OR2   \PCI-AD/IO15/$1I2246/$1I8  (
    .I0(\PCI-AD/IO15/$1I2246/M1 ),
    .I1(\PCI-AD/IO15/$1I2246/M0 ),
    .O(ADOUT15)
  );
  X_AND2   \PCI-AD/IO15/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/IO15/$1I2246/$1I7/I0 ),
    .I1(\PCI-AD/D_SLO15 ),
    .O(\PCI-AD/IO15/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD/IO4/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT4),
    .O(AD_O4),
    .RST(GND)
  );
  X_AND2   \PCI-AD/IO4/$1I2246/$1I9  (
    .I0(FAIL_ADH36),
    .I1(FAIL64_INT),
    .O(\PCI-AD/IO4/$1I2246/M1 )
  );
  X_OR2   \PCI-AD/IO4/$1I2246/$1I8  (
    .I0(\PCI-AD/IO4/$1I2246/M1 ),
    .I1(\PCI-AD/IO4/$1I2246/M0 ),
    .O(ADOUT4)
  );
  X_AND2   \PCI-AD/IO4/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/IO4/$1I2246/$1I7/I0 ),
    .I1(\PCI-AD/D_SLO4 ),
    .O(\PCI-AD/IO4/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD/IO6/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT6),
    .O(AD_O6),
    .RST(GND)
  );
  X_AND2   \PCI-AD/IO6/$1I2246/$1I9  (
    .I0(FAIL_ADH38),
    .I1(FAIL64_INT),
    .O(\PCI-AD/IO6/$1I2246/M1 )
  );
  X_OR2   \PCI-AD/IO6/$1I2246/$1I8  (
    .I0(\PCI-AD/IO6/$1I2246/M1 ),
    .I1(\PCI-AD/IO6/$1I2246/M0 ),
    .O(ADOUT6)
  );
  X_AND2   \PCI-AD/IO6/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/IO6/$1I2246/$1I7/I0 ),
    .I1(\PCI-AD/D_SLO6 ),
    .O(\PCI-AD/IO6/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD/IO5/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT5),
    .O(AD_O5),
    .RST(GND)
  );
  X_AND2   \PCI-AD/IO5/$1I2246/$1I9  (
    .I0(FAIL_ADH37),
    .I1(FAIL64_INT),
    .O(\PCI-AD/IO5/$1I2246/M1 )
  );
  X_OR2   \PCI-AD/IO5/$1I2246/$1I8  (
    .I0(\PCI-AD/IO5/$1I2246/M1 ),
    .I1(\PCI-AD/IO5/$1I2246/M0 ),
    .O(ADOUT5)
  );
  X_AND2   \PCI-AD/IO5/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/IO5/$1I2246/$1I7/I0 ),
    .I1(\PCI-AD/D_SLO5 ),
    .O(\PCI-AD/IO5/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD/IO7/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT7),
    .O(AD_O7),
    .RST(GND)
  );
  X_AND2   \PCI-AD/IO7/$1I2246/$1I9  (
    .I0(FAIL_ADH39),
    .I1(FAIL64_INT),
    .O(\PCI-AD/IO7/$1I2246/M1 )
  );
  X_OR2   \PCI-AD/IO7/$1I2246/$1I8  (
    .I0(\PCI-AD/IO7/$1I2246/M1 ),
    .I1(\PCI-AD/IO7/$1I2246/M0 ),
    .O(ADOUT7)
  );
  X_AND2   \PCI-AD/IO7/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/IO7/$1I2246/$1I7/I0 ),
    .I1(\PCI-AD/D_SLO7 ),
    .O(\PCI-AD/IO7/$1I2246/M0 )
  );
  X_AND2   \PCI-AD/$1I2927/$1I9  (
    .I0(SHADOW31),
    .I1(OUT_SEL),
    .O(\PCI-AD/$1I2927/M1 )
  );
  X_OR2   \PCI-AD/$1I2927/$1I8  (
    .I0(\PCI-AD/$1I2927/M1 ),
    .I1(\PCI-AD/$1I2927/M0 ),
    .O(\PCI-AD/D_SLO31 )
  );
  X_AND2   \PCI-AD/$1I2927/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/$1I2927/$1I7/I0 ),
    .I1(ADIO31),
    .O(\PCI-AD/$1I2927/M0 )
  );
  X_AND2   \PCI-AD/$1I2928/$1I9  (
    .I0(SHADOW30),
    .I1(OUT_SEL),
    .O(\PCI-AD/$1I2928/M1 )
  );
  X_OR2   \PCI-AD/$1I2928/$1I8  (
    .I0(\PCI-AD/$1I2928/M1 ),
    .I1(\PCI-AD/$1I2928/M0 ),
    .O(\PCI-AD/D_SLO30 )
  );
  X_AND2   \PCI-AD/$1I2928/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/$1I2928/$1I7/I0 ),
    .I1(ADIO30),
    .O(\PCI-AD/$1I2928/M0 )
  );
  X_AND2   \PCI-AD/$1I2929/$1I9  (
    .I0(SHADOW29),
    .I1(OUT_SEL),
    .O(\PCI-AD/$1I2929/M1 )
  );
  X_OR2   \PCI-AD/$1I2929/$1I8  (
    .I0(\PCI-AD/$1I2929/M1 ),
    .I1(\PCI-AD/$1I2929/M0 ),
    .O(\PCI-AD/D_SLO29 )
  );
  X_AND2   \PCI-AD/$1I2929/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/$1I2929/$1I7/I0 ),
    .I1(ADIO29),
    .O(\PCI-AD/$1I2929/M0 )
  );
  X_AND2   \PCI-AD/$1I2930/$1I9  (
    .I0(SHADOW28),
    .I1(OUT_SEL),
    .O(\PCI-AD/$1I2930/M1 )
  );
  X_OR2   \PCI-AD/$1I2930/$1I8  (
    .I0(\PCI-AD/$1I2930/M1 ),
    .I1(\PCI-AD/$1I2930/M0 ),
    .O(\PCI-AD/D_SLO28 )
  );
  X_AND2   \PCI-AD/$1I2930/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/$1I2930/$1I7/I0 ),
    .I1(ADIO28),
    .O(\PCI-AD/$1I2930/M0 )
  );
  X_AND2   \PCI-AD/$1I2931/$1I9  (
    .I0(SHADOW27),
    .I1(OUT_SEL),
    .O(\PCI-AD/$1I2931/M1 )
  );
  X_OR2   \PCI-AD/$1I2931/$1I8  (
    .I0(\PCI-AD/$1I2931/M1 ),
    .I1(\PCI-AD/$1I2931/M0 ),
    .O(\PCI-AD/D_SLO27 )
  );
  X_AND2   \PCI-AD/$1I2931/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/$1I2931/$1I7/I0 ),
    .I1(ADIO27),
    .O(\PCI-AD/$1I2931/M0 )
  );
  X_AND2   \PCI-AD/$1I2932/$1I9  (
    .I0(SHADOW26),
    .I1(OUT_SEL),
    .O(\PCI-AD/$1I2932/M1 )
  );
  X_OR2   \PCI-AD/$1I2932/$1I8  (
    .I0(\PCI-AD/$1I2932/M1 ),
    .I1(\PCI-AD/$1I2932/M0 ),
    .O(\PCI-AD/D_SLO26 )
  );
  X_AND2   \PCI-AD/$1I2932/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/$1I2932/$1I7/I0 ),
    .I1(ADIO26),
    .O(\PCI-AD/$1I2932/M0 )
  );
  X_AND2   \PCI-AD/$1I2933/$1I9  (
    .I0(SHADOW25),
    .I1(OUT_SEL),
    .O(\PCI-AD/$1I2933/M1 )
  );
  X_OR2   \PCI-AD/$1I2933/$1I8  (
    .I0(\PCI-AD/$1I2933/M1 ),
    .I1(\PCI-AD/$1I2933/M0 ),
    .O(\PCI-AD/D_SLO25 )
  );
  X_AND2   \PCI-AD/$1I2933/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/$1I2933/$1I7/I0 ),
    .I1(ADIO25),
    .O(\PCI-AD/$1I2933/M0 )
  );
  X_AND2   \PCI-AD/$1I2934/$1I9  (
    .I0(SHADOW24),
    .I1(OUT_SEL),
    .O(\PCI-AD/$1I2934/M1 )
  );
  X_OR2   \PCI-AD/$1I2934/$1I8  (
    .I0(\PCI-AD/$1I2934/M1 ),
    .I1(\PCI-AD/$1I2934/M0 ),
    .O(\PCI-AD/D_SLO24 )
  );
  X_AND2   \PCI-AD/$1I2934/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/$1I2934/$1I7/I0 ),
    .I1(ADIO24),
    .O(\PCI-AD/$1I2934/M0 )
  );
  X_AND2   \PCI-AD/$1I2935/$1I9  (
    .I0(SHADOW23),
    .I1(OUT_SEL),
    .O(\PCI-AD/$1I2935/M1 )
  );
  X_OR2   \PCI-AD/$1I2935/$1I8  (
    .I0(\PCI-AD/$1I2935/M1 ),
    .I1(\PCI-AD/$1I2935/M0 ),
    .O(\PCI-AD/D_SLO23 )
  );
  X_AND2   \PCI-AD/$1I2935/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/$1I2935/$1I7/I0 ),
    .I1(ADIO23),
    .O(\PCI-AD/$1I2935/M0 )
  );
  X_AND2   \PCI-AD/$1I2936/$1I9  (
    .I0(SHADOW22),
    .I1(OUT_SEL),
    .O(\PCI-AD/$1I2936/M1 )
  );
  X_OR2   \PCI-AD/$1I2936/$1I8  (
    .I0(\PCI-AD/$1I2936/M1 ),
    .I1(\PCI-AD/$1I2936/M0 ),
    .O(\PCI-AD/D_SLO22 )
  );
  X_AND2   \PCI-AD/$1I2936/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/$1I2936/$1I7/I0 ),
    .I1(ADIO22),
    .O(\PCI-AD/$1I2936/M0 )
  );
  X_AND2   \PCI-AD/$1I2937/$1I9  (
    .I0(SHADOW21),
    .I1(OUT_SEL),
    .O(\PCI-AD/$1I2937/M1 )
  );
  X_OR2   \PCI-AD/$1I2937/$1I8  (
    .I0(\PCI-AD/$1I2937/M1 ),
    .I1(\PCI-AD/$1I2937/M0 ),
    .O(\PCI-AD/D_SLO21 )
  );
  X_AND2   \PCI-AD/$1I2937/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/$1I2937/$1I7/I0 ),
    .I1(ADIO21),
    .O(\PCI-AD/$1I2937/M0 )
  );
  X_AND2   \PCI-AD/$1I2938/$1I9  (
    .I0(SHADOW20),
    .I1(OUT_SEL),
    .O(\PCI-AD/$1I2938/M1 )
  );
  X_OR2   \PCI-AD/$1I2938/$1I8  (
    .I0(\PCI-AD/$1I2938/M1 ),
    .I1(\PCI-AD/$1I2938/M0 ),
    .O(\PCI-AD/D_SLO20 )
  );
  X_AND2   \PCI-AD/$1I2938/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/$1I2938/$1I7/I0 ),
    .I1(ADIO20),
    .O(\PCI-AD/$1I2938/M0 )
  );
  X_AND2   \PCI-AD/$1I2939/$1I9  (
    .I0(SHADOW19),
    .I1(OUT_SEL),
    .O(\PCI-AD/$1I2939/M1 )
  );
  X_OR2   \PCI-AD/$1I2939/$1I8  (
    .I0(\PCI-AD/$1I2939/M1 ),
    .I1(\PCI-AD/$1I2939/M0 ),
    .O(\PCI-AD/D_SLO19 )
  );
  X_AND2   \PCI-AD/$1I2939/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/$1I2939/$1I7/I0 ),
    .I1(ADIO19),
    .O(\PCI-AD/$1I2939/M0 )
  );
  X_AND2   \PCI-AD/$1I2940/$1I9  (
    .I0(SHADOW18),
    .I1(OUT_SEL),
    .O(\PCI-AD/$1I2940/M1 )
  );
  X_OR2   \PCI-AD/$1I2940/$1I8  (
    .I0(\PCI-AD/$1I2940/M1 ),
    .I1(\PCI-AD/$1I2940/M0 ),
    .O(\PCI-AD/D_SLO18 )
  );
  X_AND2   \PCI-AD/$1I2940/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/$1I2940/$1I7/I0 ),
    .I1(ADIO18),
    .O(\PCI-AD/$1I2940/M0 )
  );
  X_AND2   \PCI-AD/$1I2941/$1I9  (
    .I0(SHADOW17),
    .I1(OUT_SEL),
    .O(\PCI-AD/$1I2941/M1 )
  );
  X_OR2   \PCI-AD/$1I2941/$1I8  (
    .I0(\PCI-AD/$1I2941/M1 ),
    .I1(\PCI-AD/$1I2941/M0 ),
    .O(\PCI-AD/D_SLO17 )
  );
  X_AND2   \PCI-AD/$1I2941/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/$1I2941/$1I7/I0 ),
    .I1(ADIO17),
    .O(\PCI-AD/$1I2941/M0 )
  );
  X_AND2   \PCI-AD/$1I2942/$1I9  (
    .I0(SHADOW16),
    .I1(OUT_SEL),
    .O(\PCI-AD/$1I2942/M1 )
  );
  X_OR2   \PCI-AD/$1I2942/$1I8  (
    .I0(\PCI-AD/$1I2942/M1 ),
    .I1(\PCI-AD/$1I2942/M0 ),
    .O(\PCI-AD/D_SLO16 )
  );
  X_AND2   \PCI-AD/$1I2942/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/$1I2942/$1I7/I0 ),
    .I1(ADIO16),
    .O(\PCI-AD/$1I2942/M0 )
  );
  X_AND2   \PCI-AD/$1I2943/$1I9  (
    .I0(SHADOW15),
    .I1(OUT_SEL),
    .O(\PCI-AD/$1I2943/M1 )
  );
  X_OR2   \PCI-AD/$1I2943/$1I8  (
    .I0(\PCI-AD/$1I2943/M1 ),
    .I1(\PCI-AD/$1I2943/M0 ),
    .O(\PCI-AD/D_SLO15 )
  );
  X_AND2   \PCI-AD/$1I2943/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/$1I2943/$1I7/I0 ),
    .I1(ADIO15),
    .O(\PCI-AD/$1I2943/M0 )
  );
  X_AND2   \PCI-AD/$1I2944/$1I9  (
    .I0(SHADOW14),
    .I1(OUT_SEL),
    .O(\PCI-AD/$1I2944/M1 )
  );
  X_OR2   \PCI-AD/$1I2944/$1I8  (
    .I0(\PCI-AD/$1I2944/M1 ),
    .I1(\PCI-AD/$1I2944/M0 ),
    .O(\PCI-AD/D_SLO14 )
  );
  X_AND2   \PCI-AD/$1I2944/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/$1I2944/$1I7/I0 ),
    .I1(ADIO14),
    .O(\PCI-AD/$1I2944/M0 )
  );
  X_AND2   \PCI-AD/$1I2945/$1I9  (
    .I0(SHADOW13),
    .I1(OUT_SEL),
    .O(\PCI-AD/$1I2945/M1 )
  );
  X_OR2   \PCI-AD/$1I2945/$1I8  (
    .I0(\PCI-AD/$1I2945/M1 ),
    .I1(\PCI-AD/$1I2945/M0 ),
    .O(\PCI-AD/D_SLO13 )
  );
  X_AND2   \PCI-AD/$1I2945/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/$1I2945/$1I7/I0 ),
    .I1(ADIO13),
    .O(\PCI-AD/$1I2945/M0 )
  );
  X_AND2   \PCI-AD/$1I2946/$1I9  (
    .I0(SHADOW12),
    .I1(OUT_SEL),
    .O(\PCI-AD/$1I2946/M1 )
  );
  X_OR2   \PCI-AD/$1I2946/$1I8  (
    .I0(\PCI-AD/$1I2946/M1 ),
    .I1(\PCI-AD/$1I2946/M0 ),
    .O(\PCI-AD/D_SLO12 )
  );
  X_AND2   \PCI-AD/$1I2946/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/$1I2946/$1I7/I0 ),
    .I1(ADIO12),
    .O(\PCI-AD/$1I2946/M0 )
  );
  X_AND2   \PCI-AD/$1I2947/$1I9  (
    .I0(SHADOW11),
    .I1(OUT_SEL),
    .O(\PCI-AD/$1I2947/M1 )
  );
  X_OR2   \PCI-AD/$1I2947/$1I8  (
    .I0(\PCI-AD/$1I2947/M1 ),
    .I1(\PCI-AD/$1I2947/M0 ),
    .O(\PCI-AD/D_SLO11 )
  );
  X_AND2   \PCI-AD/$1I2947/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/$1I2947/$1I7/I0 ),
    .I1(ADIO11),
    .O(\PCI-AD/$1I2947/M0 )
  );
  X_AND2   \PCI-AD/$1I2948/$1I9  (
    .I0(SHADOW10),
    .I1(OUT_SEL),
    .O(\PCI-AD/$1I2948/M1 )
  );
  X_OR2   \PCI-AD/$1I2948/$1I8  (
    .I0(\PCI-AD/$1I2948/M1 ),
    .I1(\PCI-AD/$1I2948/M0 ),
    .O(\PCI-AD/D_SLO10 )
  );
  X_AND2   \PCI-AD/$1I2948/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/$1I2948/$1I7/I0 ),
    .I1(ADIO10),
    .O(\PCI-AD/$1I2948/M0 )
  );
  X_AND2   \PCI-AD/$1I2949/$1I9  (
    .I0(SHADOW9),
    .I1(OUT_SEL),
    .O(\PCI-AD/$1I2949/M1 )
  );
  X_OR2   \PCI-AD/$1I2949/$1I8  (
    .I0(\PCI-AD/$1I2949/M1 ),
    .I1(\PCI-AD/$1I2949/M0 ),
    .O(\PCI-AD/D_SLO9 )
  );
  X_AND2   \PCI-AD/$1I2949/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/$1I2949/$1I7/I0 ),
    .I1(ADIO9),
    .O(\PCI-AD/$1I2949/M0 )
  );
  X_AND2   \PCI-AD/$1I2950/$1I9  (
    .I0(SHADOW8),
    .I1(OUT_SEL),
    .O(\PCI-AD/$1I2950/M1 )
  );
  X_OR2   \PCI-AD/$1I2950/$1I8  (
    .I0(\PCI-AD/$1I2950/M1 ),
    .I1(\PCI-AD/$1I2950/M0 ),
    .O(\PCI-AD/D_SLO8 )
  );
  X_AND2   \PCI-AD/$1I2950/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/$1I2950/$1I7/I0 ),
    .I1(ADIO8),
    .O(\PCI-AD/$1I2950/M0 )
  );
  X_AND2   \PCI-AD/$1I2951/$1I9  (
    .I0(SHADOW7),
    .I1(OUT_SEL),
    .O(\PCI-AD/$1I2951/M1 )
  );
  X_OR2   \PCI-AD/$1I2951/$1I8  (
    .I0(\PCI-AD/$1I2951/M1 ),
    .I1(\PCI-AD/$1I2951/M0 ),
    .O(\PCI-AD/D_SLO7 )
  );
  X_AND2   \PCI-AD/$1I2951/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/$1I2951/$1I7/I0 ),
    .I1(ADIO7),
    .O(\PCI-AD/$1I2951/M0 )
  );
  X_AND2   \PCI-AD/$1I2952/$1I9  (
    .I0(SHADOW6),
    .I1(OUT_SEL),
    .O(\PCI-AD/$1I2952/M1 )
  );
  X_OR2   \PCI-AD/$1I2952/$1I8  (
    .I0(\PCI-AD/$1I2952/M1 ),
    .I1(\PCI-AD/$1I2952/M0 ),
    .O(\PCI-AD/D_SLO6 )
  );
  X_AND2   \PCI-AD/$1I2952/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/$1I2952/$1I7/I0 ),
    .I1(ADIO6),
    .O(\PCI-AD/$1I2952/M0 )
  );
  X_AND2   \PCI-AD/$1I2953/$1I9  (
    .I0(SHADOW5),
    .I1(OUT_SEL),
    .O(\PCI-AD/$1I2953/M1 )
  );
  X_OR2   \PCI-AD/$1I2953/$1I8  (
    .I0(\PCI-AD/$1I2953/M1 ),
    .I1(\PCI-AD/$1I2953/M0 ),
    .O(\PCI-AD/D_SLO5 )
  );
  X_AND2   \PCI-AD/$1I2953/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/$1I2953/$1I7/I0 ),
    .I1(ADIO5),
    .O(\PCI-AD/$1I2953/M0 )
  );
  X_AND2   \PCI-AD/$1I2954/$1I9  (
    .I0(SHADOW4),
    .I1(OUT_SEL),
    .O(\PCI-AD/$1I2954/M1 )
  );
  X_OR2   \PCI-AD/$1I2954/$1I8  (
    .I0(\PCI-AD/$1I2954/M1 ),
    .I1(\PCI-AD/$1I2954/M0 ),
    .O(\PCI-AD/D_SLO4 )
  );
  X_AND2   \PCI-AD/$1I2954/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/$1I2954/$1I7/I0 ),
    .I1(ADIO4),
    .O(\PCI-AD/$1I2954/M0 )
  );
  X_AND2   \PCI-AD/$1I2955/$1I9  (
    .I0(SHADOW3),
    .I1(OUT_SEL),
    .O(\PCI-AD/$1I2955/M1 )
  );
  X_OR2   \PCI-AD/$1I2955/$1I8  (
    .I0(\PCI-AD/$1I2955/M1 ),
    .I1(\PCI-AD/$1I2955/M0 ),
    .O(\PCI-AD/D_SLO3 )
  );
  X_AND2   \PCI-AD/$1I2955/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/$1I2955/$1I7/I0 ),
    .I1(ADIO3),
    .O(\PCI-AD/$1I2955/M0 )
  );
  X_AND2   \PCI-AD/$1I2956/$1I9  (
    .I0(SHADOW2),
    .I1(OUT_SEL),
    .O(\PCI-AD/$1I2956/M1 )
  );
  X_OR2   \PCI-AD/$1I2956/$1I8  (
    .I0(\PCI-AD/$1I2956/M1 ),
    .I1(\PCI-AD/$1I2956/M0 ),
    .O(\PCI-AD/D_SLO2 )
  );
  X_AND2   \PCI-AD/$1I2956/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/$1I2956/$1I7/I0 ),
    .I1(ADIO2),
    .O(\PCI-AD/$1I2956/M0 )
  );
  X_AND2   \PCI-AD/$1I2957/$1I9  (
    .I0(SHADOW1),
    .I1(OUT_SEL),
    .O(\PCI-AD/$1I2957/M1 )
  );
  X_OR2   \PCI-AD/$1I2957/$1I8  (
    .I0(\PCI-AD/$1I2957/M1 ),
    .I1(\PCI-AD/$1I2957/M0 ),
    .O(\PCI-AD/D_SLO1 )
  );
  X_AND2   \PCI-AD/$1I2957/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/$1I2957/$1I7/I0 ),
    .I1(ADIO1),
    .O(\PCI-AD/$1I2957/M0 )
  );
  X_AND2   \PCI-AD/$1I2958/$1I9  (
    .I0(SHADOW0),
    .I1(OUT_SEL),
    .O(\PCI-AD/$1I2958/M1 )
  );
  X_OR2   \PCI-AD/$1I2958/$1I8  (
    .I0(\PCI-AD/$1I2958/M1 ),
    .I1(\PCI-AD/$1I2958/M0 ),
    .O(\PCI-AD/D_SLO0 )
  );
  X_AND2   \PCI-AD/$1I2958/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/$1I2958/$1I7/I0 ),
    .I1(ADIO0),
    .O(\PCI-AD/$1I2958/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD/IO27/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT27),
    .O(AD_O27),
    .RST(GND)
  );
  X_AND2   \PCI-AD/IO27/$1I2246/$1I9  (
    .I0(FAIL_ADH59),
    .I1(FAIL64_INT),
    .O(\PCI-AD/IO27/$1I2246/M1 )
  );
  X_OR2   \PCI-AD/IO27/$1I2246/$1I8  (
    .I0(\PCI-AD/IO27/$1I2246/M1 ),
    .I1(\PCI-AD/IO27/$1I2246/M0 ),
    .O(ADOUT27)
  );
  X_AND2   \PCI-AD/IO27/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/IO27/$1I2246/$1I7/I0 ),
    .I1(\PCI-AD/D_SLO27 ),
    .O(\PCI-AD/IO27/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD/IO26/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT26),
    .O(AD_O26),
    .RST(GND)
  );
  X_AND2   \PCI-AD/IO26/$1I2246/$1I9  (
    .I0(FAIL_ADH58),
    .I1(FAIL64_INT),
    .O(\PCI-AD/IO26/$1I2246/M1 )
  );
  X_OR2   \PCI-AD/IO26/$1I2246/$1I8  (
    .I0(\PCI-AD/IO26/$1I2246/M1 ),
    .I1(\PCI-AD/IO26/$1I2246/M0 ),
    .O(ADOUT26)
  );
  X_AND2   \PCI-AD/IO26/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/IO26/$1I2246/$1I7/I0 ),
    .I1(\PCI-AD/D_SLO26 ),
    .O(\PCI-AD/IO26/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD/IO25/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT25),
    .O(AD_O25),
    .RST(GND)
  );
  X_AND2   \PCI-AD/IO25/$1I2246/$1I9  (
    .I0(FAIL_ADH57),
    .I1(FAIL64_INT),
    .O(\PCI-AD/IO25/$1I2246/M1 )
  );
  X_OR2   \PCI-AD/IO25/$1I2246/$1I8  (
    .I0(\PCI-AD/IO25/$1I2246/M1 ),
    .I1(\PCI-AD/IO25/$1I2246/M0 ),
    .O(ADOUT25)
  );
  X_AND2   \PCI-AD/IO25/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/IO25/$1I2246/$1I7/I0 ),
    .I1(\PCI-AD/D_SLO25 ),
    .O(\PCI-AD/IO25/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD/IO24/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT24),
    .O(AD_O24),
    .RST(GND)
  );
  X_AND2   \PCI-AD/IO24/$1I2246/$1I9  (
    .I0(FAIL_ADH56),
    .I1(FAIL64_INT),
    .O(\PCI-AD/IO24/$1I2246/M1 )
  );
  X_OR2   \PCI-AD/IO24/$1I2246/$1I8  (
    .I0(\PCI-AD/IO24/$1I2246/M1 ),
    .I1(\PCI-AD/IO24/$1I2246/M0 ),
    .O(ADOUT24)
  );
  X_AND2   \PCI-AD/IO24/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/IO24/$1I2246/$1I7/I0 ),
    .I1(\PCI-AD/D_SLO24 ),
    .O(\PCI-AD/IO24/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD/IO19/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT19),
    .O(AD_O19),
    .RST(GND)
  );
  X_AND2   \PCI-AD/IO19/$1I2246/$1I9  (
    .I0(FAIL_ADH51),
    .I1(FAIL64_INT),
    .O(\PCI-AD/IO19/$1I2246/M1 )
  );
  X_OR2   \PCI-AD/IO19/$1I2246/$1I8  (
    .I0(\PCI-AD/IO19/$1I2246/M1 ),
    .I1(\PCI-AD/IO19/$1I2246/M0 ),
    .O(ADOUT19)
  );
  X_AND2   \PCI-AD/IO19/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/IO19/$1I2246/$1I7/I0 ),
    .I1(\PCI-AD/D_SLO19 ),
    .O(\PCI-AD/IO19/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD/IO18/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT18),
    .O(AD_O18),
    .RST(GND)
  );
  X_AND2   \PCI-AD/IO18/$1I2246/$1I9  (
    .I0(FAIL_ADH50),
    .I1(FAIL64_INT),
    .O(\PCI-AD/IO18/$1I2246/M1 )
  );
  X_OR2   \PCI-AD/IO18/$1I2246/$1I8  (
    .I0(\PCI-AD/IO18/$1I2246/M1 ),
    .I1(\PCI-AD/IO18/$1I2246/M0 ),
    .O(ADOUT18)
  );
  X_AND2   \PCI-AD/IO18/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/IO18/$1I2246/$1I7/I0 ),
    .I1(\PCI-AD/D_SLO18 ),
    .O(\PCI-AD/IO18/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD/IO17/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT17),
    .O(AD_O17),
    .RST(GND)
  );
  X_AND2   \PCI-AD/IO17/$1I2246/$1I9  (
    .I0(FAIL_ADH49),
    .I1(FAIL64_INT),
    .O(\PCI-AD/IO17/$1I2246/M1 )
  );
  X_OR2   \PCI-AD/IO17/$1I2246/$1I8  (
    .I0(\PCI-AD/IO17/$1I2246/M1 ),
    .I1(\PCI-AD/IO17/$1I2246/M0 ),
    .O(ADOUT17)
  );
  X_AND2   \PCI-AD/IO17/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/IO17/$1I2246/$1I7/I0 ),
    .I1(\PCI-AD/D_SLO17 ),
    .O(\PCI-AD/IO17/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD/IO16/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT16),
    .O(AD_O16),
    .RST(GND)
  );
  X_AND2   \PCI-AD/IO16/$1I2246/$1I9  (
    .I0(FAIL_ADH48),
    .I1(FAIL64_INT),
    .O(\PCI-AD/IO16/$1I2246/M1 )
  );
  X_OR2   \PCI-AD/IO16/$1I2246/$1I8  (
    .I0(\PCI-AD/IO16/$1I2246/M1 ),
    .I1(\PCI-AD/IO16/$1I2246/M0 ),
    .O(ADOUT16)
  );
  X_AND2   \PCI-AD/IO16/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/IO16/$1I2246/$1I7/I0 ),
    .I1(\PCI-AD/D_SLO16 ),
    .O(\PCI-AD/IO16/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD/IO11/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT11),
    .O(AD_O11),
    .RST(GND)
  );
  X_AND2   \PCI-AD/IO11/$1I2246/$1I9  (
    .I0(FAIL_ADH43),
    .I1(FAIL64_INT),
    .O(\PCI-AD/IO11/$1I2246/M1 )
  );
  X_OR2   \PCI-AD/IO11/$1I2246/$1I8  (
    .I0(\PCI-AD/IO11/$1I2246/M1 ),
    .I1(\PCI-AD/IO11/$1I2246/M0 ),
    .O(ADOUT11)
  );
  X_AND2   \PCI-AD/IO11/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/IO11/$1I2246/$1I7/I0 ),
    .I1(\PCI-AD/D_SLO11 ),
    .O(\PCI-AD/IO11/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD/IO10/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT10),
    .O(AD_O10),
    .RST(GND)
  );
  X_AND2   \PCI-AD/IO10/$1I2246/$1I9  (
    .I0(FAIL_ADH42),
    .I1(FAIL64_INT),
    .O(\PCI-AD/IO10/$1I2246/M1 )
  );
  X_OR2   \PCI-AD/IO10/$1I2246/$1I8  (
    .I0(\PCI-AD/IO10/$1I2246/M1 ),
    .I1(\PCI-AD/IO10/$1I2246/M0 ),
    .O(ADOUT10)
  );
  X_AND2   \PCI-AD/IO10/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/IO10/$1I2246/$1I7/I0 ),
    .I1(\PCI-AD/D_SLO10 ),
    .O(\PCI-AD/IO10/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD/IO9/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT9),
    .O(AD_O9),
    .RST(GND)
  );
  X_AND2   \PCI-AD/IO9/$1I2246/$1I9  (
    .I0(FAIL_ADH41),
    .I1(FAIL64_INT),
    .O(\PCI-AD/IO9/$1I2246/M1 )
  );
  X_OR2   \PCI-AD/IO9/$1I2246/$1I8  (
    .I0(\PCI-AD/IO9/$1I2246/M1 ),
    .I1(\PCI-AD/IO9/$1I2246/M0 ),
    .O(ADOUT9)
  );
  X_AND2   \PCI-AD/IO9/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/IO9/$1I2246/$1I7/I0 ),
    .I1(\PCI-AD/D_SLO9 ),
    .O(\PCI-AD/IO9/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD/IO8/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT8),
    .O(AD_O8),
    .RST(GND)
  );
  X_AND2   \PCI-AD/IO8/$1I2246/$1I9  (
    .I0(FAIL_ADH40),
    .I1(FAIL64_INT),
    .O(\PCI-AD/IO8/$1I2246/M1 )
  );
  X_OR2   \PCI-AD/IO8/$1I2246/$1I8  (
    .I0(\PCI-AD/IO8/$1I2246/M1 ),
    .I1(\PCI-AD/IO8/$1I2246/M0 ),
    .O(ADOUT8)
  );
  X_AND2   \PCI-AD/IO8/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/IO8/$1I2246/$1I7/I0 ),
    .I1(\PCI-AD/D_SLO8 ),
    .O(\PCI-AD/IO8/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD/IO3/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT3),
    .O(AD_O3),
    .RST(GND)
  );
  X_AND2   \PCI-AD/IO3/$1I2246/$1I9  (
    .I0(FAIL_ADH35),
    .I1(FAIL64_INT),
    .O(\PCI-AD/IO3/$1I2246/M1 )
  );
  X_OR2   \PCI-AD/IO3/$1I2246/$1I8  (
    .I0(\PCI-AD/IO3/$1I2246/M1 ),
    .I1(\PCI-AD/IO3/$1I2246/M0 ),
    .O(ADOUT3)
  );
  X_AND2   \PCI-AD/IO3/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/IO3/$1I2246/$1I7/I0 ),
    .I1(\PCI-AD/D_SLO3 ),
    .O(\PCI-AD/IO3/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD/IO2/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT2),
    .O(AD_O2),
    .RST(GND)
  );
  X_AND2   \PCI-AD/IO2/$1I2246/$1I9  (
    .I0(FAIL_ADH34),
    .I1(FAIL64_INT),
    .O(\PCI-AD/IO2/$1I2246/M1 )
  );
  X_OR2   \PCI-AD/IO2/$1I2246/$1I8  (
    .I0(\PCI-AD/IO2/$1I2246/M1 ),
    .I1(\PCI-AD/IO2/$1I2246/M0 ),
    .O(ADOUT2)
  );
  X_AND2   \PCI-AD/IO2/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/IO2/$1I2246/$1I7/I0 ),
    .I1(\PCI-AD/D_SLO2 ),
    .O(\PCI-AD/IO2/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD/IO1/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT1),
    .O(AD_O1),
    .RST(GND)
  );
  X_AND2   \PCI-AD/IO1/$1I2246/$1I9  (
    .I0(FAIL_ADH33),
    .I1(FAIL64_INT),
    .O(\PCI-AD/IO1/$1I2246/M1 )
  );
  X_OR2   \PCI-AD/IO1/$1I2246/$1I8  (
    .I0(\PCI-AD/IO1/$1I2246/M1 ),
    .I1(\PCI-AD/IO1/$1I2246/M0 ),
    .O(ADOUT1)
  );
  X_AND2   \PCI-AD/IO1/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/IO1/$1I2246/$1I7/I0 ),
    .I1(\PCI-AD/D_SLO1 ),
    .O(\PCI-AD/IO1/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD/IO0/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT0),
    .O(AD_O0),
    .RST(GND)
  );
  X_AND2   \PCI-AD/IO0/$1I2246/$1I9  (
    .I0(FAIL_ADH32),
    .I1(FAIL64_INT),
    .O(\PCI-AD/IO0/$1I2246/M1 )
  );
  X_OR2   \PCI-AD/IO0/$1I2246/$1I8  (
    .I0(\PCI-AD/IO0/$1I2246/M1 ),
    .I1(\PCI-AD/IO0/$1I2246/M0 ),
    .O(ADOUT0)
  );
  X_AND2   \PCI-AD/IO0/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD/IO0/$1I2246/$1I7/I0 ),
    .I1(\PCI-AD/D_SLO0 ),
    .O(\PCI-AD/IO0/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD_CBE/Q1  (
    .CE(SHADOW_CE),
    .CLK(CLK),
    .I(M_CBE_INT1),
    .O(SHADOW_CBE1),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD_CBE/Q3  (
    .CE(SHADOW_CE),
    .CLK(CLK),
    .I(M_CBE_INT3),
    .O(SHADOW_CBE3),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD_CBE/Q0  (
    .CE(SHADOW_CE),
    .CLK(CLK),
    .I(M_CBE_INT0),
    .O(SHADOW_CBE0),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD_CBE/Q2  (
    .CE(SHADOW_CE),
    .CLK(CLK),
    .I(M_CBE_INT2),
    .O(SHADOW_CBE2),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD/UPPER/Q15  (
    .CE(SHADOW_CE),
    .CLK(CLK),
    .I(ADIO31),
    .O(SHADOW31),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD/UPPER/Q9  (
    .CE(SHADOW_CE),
    .CLK(CLK),
    .I(ADIO25),
    .O(SHADOW25),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD/UPPER/Q13  (
    .CE(SHADOW_CE),
    .CLK(CLK),
    .I(ADIO29),
    .O(SHADOW29),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD/UPPER/Q10  (
    .CE(SHADOW_CE),
    .CLK(CLK),
    .I(ADIO26),
    .O(SHADOW26),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD/UPPER/Q14  (
    .CE(SHADOW_CE),
    .CLK(CLK),
    .I(ADIO30),
    .O(SHADOW30),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD/UPPER/Q12  (
    .CE(SHADOW_CE),
    .CLK(CLK),
    .I(ADIO28),
    .O(SHADOW28),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD/UPPER/Q11  (
    .CE(SHADOW_CE),
    .CLK(CLK),
    .I(ADIO27),
    .O(SHADOW27),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD/UPPER/Q8  (
    .CE(SHADOW_CE),
    .CLK(CLK),
    .I(ADIO24),
    .O(SHADOW24),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD/UPPER/Q7  (
    .CE(SHADOW_CE),
    .CLK(CLK),
    .I(ADIO23),
    .O(SHADOW23),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD/UPPER/Q1  (
    .CE(SHADOW_CE),
    .CLK(CLK),
    .I(ADIO17),
    .O(SHADOW17),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD/UPPER/Q5  (
    .CE(SHADOW_CE),
    .CLK(CLK),
    .I(ADIO21),
    .O(SHADOW21),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD/UPPER/Q3  (
    .CE(SHADOW_CE),
    .CLK(CLK),
    .I(ADIO19),
    .O(SHADOW19),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD/UPPER/Q0  (
    .CE(SHADOW_CE),
    .CLK(CLK),
    .I(ADIO16),
    .O(SHADOW16),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD/UPPER/Q2  (
    .CE(SHADOW_CE),
    .CLK(CLK),
    .I(ADIO18),
    .O(SHADOW18),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD/UPPER/Q4  (
    .CE(SHADOW_CE),
    .CLK(CLK),
    .I(ADIO20),
    .O(SHADOW20),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD/UPPER/Q6  (
    .CE(SHADOW_CE),
    .CLK(CLK),
    .I(ADIO22),
    .O(SHADOW22),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD/LOWER/Q15  (
    .CE(SHADOW_CE),
    .CLK(CLK),
    .I(ADIO15),
    .O(SHADOW15),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD/LOWER/Q9  (
    .CE(SHADOW_CE),
    .CLK(CLK),
    .I(ADIO9),
    .O(SHADOW9),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD/LOWER/Q13  (
    .CE(SHADOW_CE),
    .CLK(CLK),
    .I(ADIO13),
    .O(SHADOW13),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD/LOWER/Q10  (
    .CE(SHADOW_CE),
    .CLK(CLK),
    .I(ADIO10),
    .O(SHADOW10),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD/LOWER/Q14  (
    .CE(SHADOW_CE),
    .CLK(CLK),
    .I(ADIO14),
    .O(SHADOW14),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD/LOWER/Q12  (
    .CE(SHADOW_CE),
    .CLK(CLK),
    .I(ADIO12),
    .O(SHADOW12),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD/LOWER/Q11  (
    .CE(SHADOW_CE),
    .CLK(CLK),
    .I(ADIO11),
    .O(SHADOW11),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD/LOWER/Q8  (
    .CE(SHADOW_CE),
    .CLK(CLK),
    .I(ADIO8),
    .O(SHADOW8),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD/LOWER/Q7  (
    .CE(SHADOW_CE),
    .CLK(CLK),
    .I(ADIO7),
    .O(SHADOW7),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD/LOWER/Q1  (
    .CE(SHADOW_CE),
    .CLK(CLK),
    .I(ADIO1),
    .O(SHADOW1),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD/LOWER/Q5  (
    .CE(SHADOW_CE),
    .CLK(CLK),
    .I(ADIO5),
    .O(SHADOW5),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD/LOWER/Q3  (
    .CE(SHADOW_CE),
    .CLK(CLK),
    .I(ADIO3),
    .O(SHADOW3),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD/LOWER/Q0  (
    .CE(SHADOW_CE),
    .CLK(CLK),
    .I(ADIO0),
    .O(SHADOW0),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD/LOWER/Q2  (
    .CE(SHADOW_CE),
    .CLK(CLK),
    .I(ADIO2),
    .O(SHADOW2),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD/LOWER/Q4  (
    .CE(SHADOW_CE),
    .CLK(CLK),
    .I(ADIO4),
    .O(SHADOW4),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD/LOWER/Q6  (
    .CE(SHADOW_CE),
    .CLK(CLK),
    .I(ADIO6),
    .O(SHADOW6),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD64/IO28/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT60),
    .O(AD_O60),
    .RST(GND)
  );
  X_AND2   \PCI-AD64/IO28/$1I2246/$1I9  (
    .I0(SHADOW60),
    .I1(OUT_SEL64),
    .O(\PCI-AD64/IO28/$1I2246/M1 )
  );
  X_OR2   \PCI-AD64/IO28/$1I2246/$1I8  (
    .I0(\PCI-AD64/IO28/$1I2246/M1 ),
    .I1(\PCI-AD64/IO28/$1I2246/M0 ),
    .O(ADOUT60)
  );
  X_AND2   \PCI-AD64/IO28/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD64/IO28/$1I2246/$1I7/I0 ),
    .I1(ADIO60),
    .O(\PCI-AD64/IO28/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD64/IO30/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT62),
    .O(AD_O62),
    .RST(GND)
  );
  X_AND2   \PCI-AD64/IO30/$1I2246/$1I9  (
    .I0(SHADOW62),
    .I1(OUT_SEL64),
    .O(\PCI-AD64/IO30/$1I2246/M1 )
  );
  X_OR2   \PCI-AD64/IO30/$1I2246/$1I8  (
    .I0(\PCI-AD64/IO30/$1I2246/M1 ),
    .I1(\PCI-AD64/IO30/$1I2246/M0 ),
    .O(ADOUT62)
  );
  X_AND2   \PCI-AD64/IO30/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD64/IO30/$1I2246/$1I7/I0 ),
    .I1(ADIO62),
    .O(\PCI-AD64/IO30/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD64/IO29/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT61),
    .O(AD_O61),
    .RST(GND)
  );
  X_AND2   \PCI-AD64/IO29/$1I2246/$1I9  (
    .I0(SHADOW61),
    .I1(OUT_SEL64),
    .O(\PCI-AD64/IO29/$1I2246/M1 )
  );
  X_OR2   \PCI-AD64/IO29/$1I2246/$1I8  (
    .I0(\PCI-AD64/IO29/$1I2246/M1 ),
    .I1(\PCI-AD64/IO29/$1I2246/M0 ),
    .O(ADOUT61)
  );
  X_AND2   \PCI-AD64/IO29/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD64/IO29/$1I2246/$1I7/I0 ),
    .I1(ADIO61),
    .O(\PCI-AD64/IO29/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD64/IO31/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT63),
    .O(AD_O63),
    .RST(GND)
  );
  X_AND2   \PCI-AD64/IO31/$1I2246/$1I9  (
    .I0(SHADOW63),
    .I1(OUT_SEL64),
    .O(\PCI-AD64/IO31/$1I2246/M1 )
  );
  X_OR2   \PCI-AD64/IO31/$1I2246/$1I8  (
    .I0(\PCI-AD64/IO31/$1I2246/M1 ),
    .I1(\PCI-AD64/IO31/$1I2246/M0 ),
    .O(ADOUT63)
  );
  X_AND2   \PCI-AD64/IO31/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD64/IO31/$1I2246/$1I7/I0 ),
    .I1(ADIO63),
    .O(\PCI-AD64/IO31/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD64/IO20/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT52),
    .O(AD_O52),
    .RST(GND)
  );
  X_AND2   \PCI-AD64/IO20/$1I2246/$1I9  (
    .I0(SHADOW52),
    .I1(OUT_SEL64),
    .O(\PCI-AD64/IO20/$1I2246/M1 )
  );
  X_OR2   \PCI-AD64/IO20/$1I2246/$1I8  (
    .I0(\PCI-AD64/IO20/$1I2246/M1 ),
    .I1(\PCI-AD64/IO20/$1I2246/M0 ),
    .O(ADOUT52)
  );
  X_AND2   \PCI-AD64/IO20/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD64/IO20/$1I2246/$1I7/I0 ),
    .I1(ADIO52),
    .O(\PCI-AD64/IO20/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD64/IO22/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT54),
    .O(AD_O54),
    .RST(GND)
  );
  X_AND2   \PCI-AD64/IO22/$1I2246/$1I9  (
    .I0(SHADOW54),
    .I1(OUT_SEL64),
    .O(\PCI-AD64/IO22/$1I2246/M1 )
  );
  X_OR2   \PCI-AD64/IO22/$1I2246/$1I8  (
    .I0(\PCI-AD64/IO22/$1I2246/M1 ),
    .I1(\PCI-AD64/IO22/$1I2246/M0 ),
    .O(ADOUT54)
  );
  X_AND2   \PCI-AD64/IO22/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD64/IO22/$1I2246/$1I7/I0 ),
    .I1(ADIO54),
    .O(\PCI-AD64/IO22/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD64/IO21/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT53),
    .O(AD_O53),
    .RST(GND)
  );
  X_AND2   \PCI-AD64/IO21/$1I2246/$1I9  (
    .I0(SHADOW53),
    .I1(OUT_SEL64),
    .O(\PCI-AD64/IO21/$1I2246/M1 )
  );
  X_OR2   \PCI-AD64/IO21/$1I2246/$1I8  (
    .I0(\PCI-AD64/IO21/$1I2246/M1 ),
    .I1(\PCI-AD64/IO21/$1I2246/M0 ),
    .O(ADOUT53)
  );
  X_AND2   \PCI-AD64/IO21/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD64/IO21/$1I2246/$1I7/I0 ),
    .I1(ADIO53),
    .O(\PCI-AD64/IO21/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD64/IO23/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT55),
    .O(AD_O55),
    .RST(GND)
  );
  X_AND2   \PCI-AD64/IO23/$1I2246/$1I9  (
    .I0(SHADOW55),
    .I1(OUT_SEL64),
    .O(\PCI-AD64/IO23/$1I2246/M1 )
  );
  X_OR2   \PCI-AD64/IO23/$1I2246/$1I8  (
    .I0(\PCI-AD64/IO23/$1I2246/M1 ),
    .I1(\PCI-AD64/IO23/$1I2246/M0 ),
    .O(ADOUT55)
  );
  X_AND2   \PCI-AD64/IO23/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD64/IO23/$1I2246/$1I7/I0 ),
    .I1(ADIO55),
    .O(\PCI-AD64/IO23/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD64/IO12/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT44),
    .O(AD_O44),
    .RST(GND)
  );
  X_AND2   \PCI-AD64/IO12/$1I2246/$1I9  (
    .I0(SHADOW44),
    .I1(OUT_SEL64),
    .O(\PCI-AD64/IO12/$1I2246/M1 )
  );
  X_OR2   \PCI-AD64/IO12/$1I2246/$1I8  (
    .I0(\PCI-AD64/IO12/$1I2246/M1 ),
    .I1(\PCI-AD64/IO12/$1I2246/M0 ),
    .O(ADOUT44)
  );
  X_AND2   \PCI-AD64/IO12/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD64/IO12/$1I2246/$1I7/I0 ),
    .I1(ADIO44),
    .O(\PCI-AD64/IO12/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD64/IO14/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT46),
    .O(AD_O46),
    .RST(GND)
  );
  X_AND2   \PCI-AD64/IO14/$1I2246/$1I9  (
    .I0(SHADOW46),
    .I1(OUT_SEL64),
    .O(\PCI-AD64/IO14/$1I2246/M1 )
  );
  X_OR2   \PCI-AD64/IO14/$1I2246/$1I8  (
    .I0(\PCI-AD64/IO14/$1I2246/M1 ),
    .I1(\PCI-AD64/IO14/$1I2246/M0 ),
    .O(ADOUT46)
  );
  X_AND2   \PCI-AD64/IO14/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD64/IO14/$1I2246/$1I7/I0 ),
    .I1(ADIO46),
    .O(\PCI-AD64/IO14/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD64/IO13/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT45),
    .O(AD_O45),
    .RST(GND)
  );
  X_AND2   \PCI-AD64/IO13/$1I2246/$1I9  (
    .I0(SHADOW45),
    .I1(OUT_SEL64),
    .O(\PCI-AD64/IO13/$1I2246/M1 )
  );
  X_OR2   \PCI-AD64/IO13/$1I2246/$1I8  (
    .I0(\PCI-AD64/IO13/$1I2246/M1 ),
    .I1(\PCI-AD64/IO13/$1I2246/M0 ),
    .O(ADOUT45)
  );
  X_AND2   \PCI-AD64/IO13/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD64/IO13/$1I2246/$1I7/I0 ),
    .I1(ADIO45),
    .O(\PCI-AD64/IO13/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD64/IO15/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT47),
    .O(AD_O47),
    .RST(GND)
  );
  X_AND2   \PCI-AD64/IO15/$1I2246/$1I9  (
    .I0(SHADOW47),
    .I1(OUT_SEL64),
    .O(\PCI-AD64/IO15/$1I2246/M1 )
  );
  X_OR2   \PCI-AD64/IO15/$1I2246/$1I8  (
    .I0(\PCI-AD64/IO15/$1I2246/M1 ),
    .I1(\PCI-AD64/IO15/$1I2246/M0 ),
    .O(ADOUT47)
  );
  X_AND2   \PCI-AD64/IO15/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD64/IO15/$1I2246/$1I7/I0 ),
    .I1(ADIO47),
    .O(\PCI-AD64/IO15/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD64/IO4/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT36),
    .O(AD_O36),
    .RST(GND)
  );
  X_AND2   \PCI-AD64/IO4/$1I2246/$1I9  (
    .I0(SHADOW36),
    .I1(OUT_SEL64),
    .O(\PCI-AD64/IO4/$1I2246/M1 )
  );
  X_OR2   \PCI-AD64/IO4/$1I2246/$1I8  (
    .I0(\PCI-AD64/IO4/$1I2246/M1 ),
    .I1(\PCI-AD64/IO4/$1I2246/M0 ),
    .O(ADOUT36)
  );
  X_AND2   \PCI-AD64/IO4/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD64/IO4/$1I2246/$1I7/I0 ),
    .I1(ADIO36),
    .O(\PCI-AD64/IO4/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD64/IO6/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT38),
    .O(AD_O38),
    .RST(GND)
  );
  X_AND2   \PCI-AD64/IO6/$1I2246/$1I9  (
    .I0(SHADOW38),
    .I1(OUT_SEL64),
    .O(\PCI-AD64/IO6/$1I2246/M1 )
  );
  X_OR2   \PCI-AD64/IO6/$1I2246/$1I8  (
    .I0(\PCI-AD64/IO6/$1I2246/M1 ),
    .I1(\PCI-AD64/IO6/$1I2246/M0 ),
    .O(ADOUT38)
  );
  X_AND2   \PCI-AD64/IO6/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD64/IO6/$1I2246/$1I7/I0 ),
    .I1(ADIO38),
    .O(\PCI-AD64/IO6/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD64/IO5/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT37),
    .O(AD_O37),
    .RST(GND)
  );
  X_AND2   \PCI-AD64/IO5/$1I2246/$1I9  (
    .I0(SHADOW37),
    .I1(OUT_SEL64),
    .O(\PCI-AD64/IO5/$1I2246/M1 )
  );
  X_OR2   \PCI-AD64/IO5/$1I2246/$1I8  (
    .I0(\PCI-AD64/IO5/$1I2246/M1 ),
    .I1(\PCI-AD64/IO5/$1I2246/M0 ),
    .O(ADOUT37)
  );
  X_AND2   \PCI-AD64/IO5/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD64/IO5/$1I2246/$1I7/I0 ),
    .I1(ADIO37),
    .O(\PCI-AD64/IO5/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD64/IO7/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT39),
    .O(AD_O39),
    .RST(GND)
  );
  X_AND2   \PCI-AD64/IO7/$1I2246/$1I9  (
    .I0(SHADOW39),
    .I1(OUT_SEL64),
    .O(\PCI-AD64/IO7/$1I2246/M1 )
  );
  X_OR2   \PCI-AD64/IO7/$1I2246/$1I8  (
    .I0(\PCI-AD64/IO7/$1I2246/M1 ),
    .I1(\PCI-AD64/IO7/$1I2246/M0 ),
    .O(ADOUT39)
  );
  X_AND2   \PCI-AD64/IO7/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD64/IO7/$1I2246/$1I7/I0 ),
    .I1(ADIO39),
    .O(\PCI-AD64/IO7/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD64/IO27/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT59),
    .O(AD_O59),
    .RST(GND)
  );
  X_AND2   \PCI-AD64/IO27/$1I2246/$1I9  (
    .I0(SHADOW59),
    .I1(OUT_SEL64),
    .O(\PCI-AD64/IO27/$1I2246/M1 )
  );
  X_OR2   \PCI-AD64/IO27/$1I2246/$1I8  (
    .I0(\PCI-AD64/IO27/$1I2246/M1 ),
    .I1(\PCI-AD64/IO27/$1I2246/M0 ),
    .O(ADOUT59)
  );
  X_AND2   \PCI-AD64/IO27/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD64/IO27/$1I2246/$1I7/I0 ),
    .I1(ADIO59),
    .O(\PCI-AD64/IO27/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD64/IO26/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT58),
    .O(AD_O58),
    .RST(GND)
  );
  X_AND2   \PCI-AD64/IO26/$1I2246/$1I9  (
    .I0(SHADOW58),
    .I1(OUT_SEL64),
    .O(\PCI-AD64/IO26/$1I2246/M1 )
  );
  X_OR2   \PCI-AD64/IO26/$1I2246/$1I8  (
    .I0(\PCI-AD64/IO26/$1I2246/M1 ),
    .I1(\PCI-AD64/IO26/$1I2246/M0 ),
    .O(ADOUT58)
  );
  X_AND2   \PCI-AD64/IO26/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD64/IO26/$1I2246/$1I7/I0 ),
    .I1(ADIO58),
    .O(\PCI-AD64/IO26/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD64/IO25/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT57),
    .O(AD_O57),
    .RST(GND)
  );
  X_AND2   \PCI-AD64/IO25/$1I2246/$1I9  (
    .I0(SHADOW57),
    .I1(OUT_SEL64),
    .O(\PCI-AD64/IO25/$1I2246/M1 )
  );
  X_OR2   \PCI-AD64/IO25/$1I2246/$1I8  (
    .I0(\PCI-AD64/IO25/$1I2246/M1 ),
    .I1(\PCI-AD64/IO25/$1I2246/M0 ),
    .O(ADOUT57)
  );
  X_AND2   \PCI-AD64/IO25/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD64/IO25/$1I2246/$1I7/I0 ),
    .I1(ADIO57),
    .O(\PCI-AD64/IO25/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD64/IO24/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT56),
    .O(AD_O56),
    .RST(GND)
  );
  X_AND2   \PCI-AD64/IO24/$1I2246/$1I9  (
    .I0(SHADOW56),
    .I1(OUT_SEL64),
    .O(\PCI-AD64/IO24/$1I2246/M1 )
  );
  X_OR2   \PCI-AD64/IO24/$1I2246/$1I8  (
    .I0(\PCI-AD64/IO24/$1I2246/M1 ),
    .I1(\PCI-AD64/IO24/$1I2246/M0 ),
    .O(ADOUT56)
  );
  X_AND2   \PCI-AD64/IO24/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD64/IO24/$1I2246/$1I7/I0 ),
    .I1(ADIO56),
    .O(\PCI-AD64/IO24/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD64/IO19/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT51),
    .O(AD_O51),
    .RST(GND)
  );
  X_AND2   \PCI-AD64/IO19/$1I2246/$1I9  (
    .I0(SHADOW51),
    .I1(OUT_SEL64),
    .O(\PCI-AD64/IO19/$1I2246/M1 )
  );
  X_OR2   \PCI-AD64/IO19/$1I2246/$1I8  (
    .I0(\PCI-AD64/IO19/$1I2246/M1 ),
    .I1(\PCI-AD64/IO19/$1I2246/M0 ),
    .O(ADOUT51)
  );
  X_AND2   \PCI-AD64/IO19/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD64/IO19/$1I2246/$1I7/I0 ),
    .I1(ADIO51),
    .O(\PCI-AD64/IO19/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD64/IO18/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT50),
    .O(AD_O50),
    .RST(GND)
  );
  X_AND2   \PCI-AD64/IO18/$1I2246/$1I9  (
    .I0(SHADOW50),
    .I1(OUT_SEL64),
    .O(\PCI-AD64/IO18/$1I2246/M1 )
  );
  X_OR2   \PCI-AD64/IO18/$1I2246/$1I8  (
    .I0(\PCI-AD64/IO18/$1I2246/M1 ),
    .I1(\PCI-AD64/IO18/$1I2246/M0 ),
    .O(ADOUT50)
  );
  X_AND2   \PCI-AD64/IO18/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD64/IO18/$1I2246/$1I7/I0 ),
    .I1(ADIO50),
    .O(\PCI-AD64/IO18/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD64/IO17/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT49),
    .O(AD_O49),
    .RST(GND)
  );
  X_AND2   \PCI-AD64/IO17/$1I2246/$1I9  (
    .I0(SHADOW49),
    .I1(OUT_SEL64),
    .O(\PCI-AD64/IO17/$1I2246/M1 )
  );
  X_OR2   \PCI-AD64/IO17/$1I2246/$1I8  (
    .I0(\PCI-AD64/IO17/$1I2246/M1 ),
    .I1(\PCI-AD64/IO17/$1I2246/M0 ),
    .O(ADOUT49)
  );
  X_AND2   \PCI-AD64/IO17/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD64/IO17/$1I2246/$1I7/I0 ),
    .I1(ADIO49),
    .O(\PCI-AD64/IO17/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD64/IO16/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT48),
    .O(AD_O48),
    .RST(GND)
  );
  X_AND2   \PCI-AD64/IO16/$1I2246/$1I9  (
    .I0(SHADOW48),
    .I1(OUT_SEL64),
    .O(\PCI-AD64/IO16/$1I2246/M1 )
  );
  X_OR2   \PCI-AD64/IO16/$1I2246/$1I8  (
    .I0(\PCI-AD64/IO16/$1I2246/M1 ),
    .I1(\PCI-AD64/IO16/$1I2246/M0 ),
    .O(ADOUT48)
  );
  X_AND2   \PCI-AD64/IO16/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD64/IO16/$1I2246/$1I7/I0 ),
    .I1(ADIO48),
    .O(\PCI-AD64/IO16/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD64/IO11/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT43),
    .O(AD_O43),
    .RST(GND)
  );
  X_AND2   \PCI-AD64/IO11/$1I2246/$1I9  (
    .I0(SHADOW43),
    .I1(OUT_SEL64),
    .O(\PCI-AD64/IO11/$1I2246/M1 )
  );
  X_OR2   \PCI-AD64/IO11/$1I2246/$1I8  (
    .I0(\PCI-AD64/IO11/$1I2246/M1 ),
    .I1(\PCI-AD64/IO11/$1I2246/M0 ),
    .O(ADOUT43)
  );
  X_AND2   \PCI-AD64/IO11/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD64/IO11/$1I2246/$1I7/I0 ),
    .I1(ADIO43),
    .O(\PCI-AD64/IO11/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD64/IO10/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT42),
    .O(AD_O42),
    .RST(GND)
  );
  X_AND2   \PCI-AD64/IO10/$1I2246/$1I9  (
    .I0(SHADOW42),
    .I1(OUT_SEL64),
    .O(\PCI-AD64/IO10/$1I2246/M1 )
  );
  X_OR2   \PCI-AD64/IO10/$1I2246/$1I8  (
    .I0(\PCI-AD64/IO10/$1I2246/M1 ),
    .I1(\PCI-AD64/IO10/$1I2246/M0 ),
    .O(ADOUT42)
  );
  X_AND2   \PCI-AD64/IO10/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD64/IO10/$1I2246/$1I7/I0 ),
    .I1(ADIO42),
    .O(\PCI-AD64/IO10/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD64/IO9/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT41),
    .O(AD_O41),
    .RST(GND)
  );
  X_AND2   \PCI-AD64/IO9/$1I2246/$1I9  (
    .I0(SHADOW41),
    .I1(OUT_SEL64),
    .O(\PCI-AD64/IO9/$1I2246/M1 )
  );
  X_OR2   \PCI-AD64/IO9/$1I2246/$1I8  (
    .I0(\PCI-AD64/IO9/$1I2246/M1 ),
    .I1(\PCI-AD64/IO9/$1I2246/M0 ),
    .O(ADOUT41)
  );
  X_AND2   \PCI-AD64/IO9/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD64/IO9/$1I2246/$1I7/I0 ),
    .I1(ADIO41),
    .O(\PCI-AD64/IO9/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD64/IO8/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT40),
    .O(AD_O40),
    .RST(GND)
  );
  X_AND2   \PCI-AD64/IO8/$1I2246/$1I9  (
    .I0(SHADOW40),
    .I1(OUT_SEL64),
    .O(\PCI-AD64/IO8/$1I2246/M1 )
  );
  X_OR2   \PCI-AD64/IO8/$1I2246/$1I8  (
    .I0(\PCI-AD64/IO8/$1I2246/M1 ),
    .I1(\PCI-AD64/IO8/$1I2246/M0 ),
    .O(ADOUT40)
  );
  X_AND2   \PCI-AD64/IO8/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD64/IO8/$1I2246/$1I7/I0 ),
    .I1(ADIO40),
    .O(\PCI-AD64/IO8/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD64/IO3/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT35),
    .O(AD_O35),
    .RST(GND)
  );
  X_AND2   \PCI-AD64/IO3/$1I2246/$1I9  (
    .I0(SHADOW35),
    .I1(OUT_SEL64),
    .O(\PCI-AD64/IO3/$1I2246/M1 )
  );
  X_OR2   \PCI-AD64/IO3/$1I2246/$1I8  (
    .I0(\PCI-AD64/IO3/$1I2246/M1 ),
    .I1(\PCI-AD64/IO3/$1I2246/M0 ),
    .O(ADOUT35)
  );
  X_AND2   \PCI-AD64/IO3/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD64/IO3/$1I2246/$1I7/I0 ),
    .I1(ADIO35),
    .O(\PCI-AD64/IO3/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD64/IO2/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT34),
    .O(AD_O34),
    .RST(GND)
  );
  X_AND2   \PCI-AD64/IO2/$1I2246/$1I9  (
    .I0(SHADOW34),
    .I1(OUT_SEL64),
    .O(\PCI-AD64/IO2/$1I2246/M1 )
  );
  X_OR2   \PCI-AD64/IO2/$1I2246/$1I8  (
    .I0(\PCI-AD64/IO2/$1I2246/M1 ),
    .I1(\PCI-AD64/IO2/$1I2246/M0 ),
    .O(ADOUT34)
  );
  X_AND2   \PCI-AD64/IO2/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD64/IO2/$1I2246/$1I7/I0 ),
    .I1(ADIO34),
    .O(\PCI-AD64/IO2/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD64/IO1/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT33),
    .O(AD_O33),
    .RST(GND)
  );
  X_AND2   \PCI-AD64/IO1/$1I2246/$1I9  (
    .I0(SHADOW33),
    .I1(OUT_SEL64),
    .O(\PCI-AD64/IO1/$1I2246/M1 )
  );
  X_OR2   \PCI-AD64/IO1/$1I2246/$1I8  (
    .I0(\PCI-AD64/IO1/$1I2246/M1 ),
    .I1(\PCI-AD64/IO1/$1I2246/M0 ),
    .O(ADOUT33)
  );
  X_AND2   \PCI-AD64/IO1/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD64/IO1/$1I2246/$1I7/I0 ),
    .I1(ADIO33),
    .O(\PCI-AD64/IO1/$1I2246/M0 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-AD64/IO0/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(ADOUT32),
    .O(AD_O32),
    .RST(GND)
  );
  X_AND2   \PCI-AD64/IO0/$1I2246/$1I9  (
    .I0(SHADOW32),
    .I1(OUT_SEL64),
    .O(\PCI-AD64/IO0/$1I2246/M1 )
  );
  X_OR2   \PCI-AD64/IO0/$1I2246/$1I8  (
    .I0(\PCI-AD64/IO0/$1I2246/M1 ),
    .I1(\PCI-AD64/IO0/$1I2246/M0 ),
    .O(ADOUT32)
  );
  X_AND2   \PCI-AD64/IO0/$1I2246/$1I7  (
    .I0(\NlwInverterSignal_PCI-AD64/IO0/$1I2246/$1I7/I0 ),
    .I1(ADIO32),
    .O(\PCI-AD64/IO0/$1I2246/M0 )
  );
  X_AND2   \PCI-CBE64/IO3/$1I2316  (
    .I0(\PCI-CBE64/$1N2797 ),
    .I1(\PCI-CBE64/$1N2801 ),
    .O(\PCI-CBE64/IO3/$1N2321 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-CBE64/IO3/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(CBEOUT7),
    .O(CBE_O7),
    .RST(GND)
  );
  X_AND2   \PCI-CBE64/IO3/$1I2296/$1I9  (
    .I0(SHADOW_CBE7),
    .I1(OUT_SEL64),
    .O(\PCI-CBE64/IO3/$1I2296/M1 )
  );
  X_OR2   \PCI-CBE64/IO3/$1I2296/$1I8  (
    .I0(\PCI-CBE64/IO3/$1I2296/M1 ),
    .I1(\PCI-CBE64/IO3/$1I2296/M0 ),
    .O(\PCI-CBE64/IO3/D_SLO )
  );
  X_AND2   \PCI-CBE64/IO3/$1I2296/$1I7  (
    .I0(\NlwInverterSignal_PCI-CBE64/IO3/$1I2296/$1I7/I0 ),
    .I1(M_CBE_INT7),
    .O(\PCI-CBE64/IO3/$1I2296/M0 )
  );
  X_AND2   \PCI-CBE64/IO3/$1I2303/$1I9  (
    .I0(\PCI-CBE64/$1N2799 ),
    .I1(\PCI-CBE64/IO3/$1N2321 ),
    .O(\PCI-CBE64/IO3/$1I2303/M1 )
  );
  X_OR2   \PCI-CBE64/IO3/$1I2303/$1I8  (
    .I0(\PCI-CBE64/IO3/$1I2303/M1 ),
    .I1(\PCI-CBE64/IO3/$1I2303/M0 ),
    .O(CBEOUT7)
  );
  X_AND2   \PCI-CBE64/IO3/$1I2303/$1I7  (
    .I0(\NlwInverterSignal_PCI-CBE64/IO3/$1I2303/$1I7/I0 ),
    .I1(\PCI-CBE64/IO3/D_SLO ),
    .O(\PCI-CBE64/IO3/$1I2303/M0 )
  );
  X_AND2   \PCI-CBE64/IO2/$1I2316  (
    .I0(\PCI-CBE64/$1N2791 ),
    .I1(\PCI-CBE64/$1N2795 ),
    .O(\PCI-CBE64/IO2/$1N2321 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-CBE64/IO2/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(CBEOUT6),
    .O(CBE_O6),
    .RST(GND)
  );
  X_AND2   \PCI-CBE64/IO2/$1I2296/$1I9  (
    .I0(SHADOW_CBE6),
    .I1(OUT_SEL64),
    .O(\PCI-CBE64/IO2/$1I2296/M1 )
  );
  X_OR2   \PCI-CBE64/IO2/$1I2296/$1I8  (
    .I0(\PCI-CBE64/IO2/$1I2296/M1 ),
    .I1(\PCI-CBE64/IO2/$1I2296/M0 ),
    .O(\PCI-CBE64/IO2/D_SLO )
  );
  X_AND2   \PCI-CBE64/IO2/$1I2296/$1I7  (
    .I0(\NlwInverterSignal_PCI-CBE64/IO2/$1I2296/$1I7/I0 ),
    .I1(M_CBE_INT6),
    .O(\PCI-CBE64/IO2/$1I2296/M0 )
  );
  X_AND2   \PCI-CBE64/IO2/$1I2303/$1I9  (
    .I0(\PCI-CBE64/$1N2793 ),
    .I1(\PCI-CBE64/IO2/$1N2321 ),
    .O(\PCI-CBE64/IO2/$1I2303/M1 )
  );
  X_OR2   \PCI-CBE64/IO2/$1I2303/$1I8  (
    .I0(\PCI-CBE64/IO2/$1I2303/M1 ),
    .I1(\PCI-CBE64/IO2/$1I2303/M0 ),
    .O(CBEOUT6)
  );
  X_AND2   \PCI-CBE64/IO2/$1I2303/$1I7  (
    .I0(\NlwInverterSignal_PCI-CBE64/IO2/$1I2303/$1I7/I0 ),
    .I1(\PCI-CBE64/IO2/D_SLO ),
    .O(\PCI-CBE64/IO2/$1I2303/M0 )
  );
  X_AND2   \PCI-CBE64/IO1/$1I2316  (
    .I0(\PCI-CBE64/$1N2785 ),
    .I1(\PCI-CBE64/$1N2789 ),
    .O(\PCI-CBE64/IO1/$1N2321 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-CBE64/IO1/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(CBEOUT5),
    .O(CBE_O5),
    .RST(GND)
  );
  X_AND2   \PCI-CBE64/IO1/$1I2296/$1I9  (
    .I0(SHADOW_CBE5),
    .I1(OUT_SEL64),
    .O(\PCI-CBE64/IO1/$1I2296/M1 )
  );
  X_OR2   \PCI-CBE64/IO1/$1I2296/$1I8  (
    .I0(\PCI-CBE64/IO1/$1I2296/M1 ),
    .I1(\PCI-CBE64/IO1/$1I2296/M0 ),
    .O(\PCI-CBE64/IO1/D_SLO )
  );
  X_AND2   \PCI-CBE64/IO1/$1I2296/$1I7  (
    .I0(\NlwInverterSignal_PCI-CBE64/IO1/$1I2296/$1I7/I0 ),
    .I1(M_CBE_INT5),
    .O(\PCI-CBE64/IO1/$1I2296/M0 )
  );
  X_AND2   \PCI-CBE64/IO1/$1I2303/$1I9  (
    .I0(\PCI-CBE64/$1N2787 ),
    .I1(\PCI-CBE64/IO1/$1N2321 ),
    .O(\PCI-CBE64/IO1/$1I2303/M1 )
  );
  X_OR2   \PCI-CBE64/IO1/$1I2303/$1I8  (
    .I0(\PCI-CBE64/IO1/$1I2303/M1 ),
    .I1(\PCI-CBE64/IO1/$1I2303/M0 ),
    .O(CBEOUT5)
  );
  X_AND2   \PCI-CBE64/IO1/$1I2303/$1I7  (
    .I0(\NlwInverterSignal_PCI-CBE64/IO1/$1I2303/$1I7/I0 ),
    .I1(\PCI-CBE64/IO1/D_SLO ),
    .O(\PCI-CBE64/IO1/$1I2303/M0 )
  );
  X_AND2   \PCI-CBE64/IO0/$1I2316  (
    .I0(\PCI-CBE64/$1N2779 ),
    .I1(\PCI-CBE64/$1N2783 ),
    .O(\PCI-CBE64/IO0/$1N2321 )
  );
  X_FF #(
    .INIT ( 1'b1 ))
  \PCI-CBE64/IO0/OFD  (
    .SET(NlwRenamedSig_OI_RST),
    .CE(PCI_CE),
    .CLK(CLKX),
    .I(CBEOUT4),
    .O(CBE_O4),
    .RST(GND)
  );
  X_AND2   \PCI-CBE64/IO0/$1I2296/$1I9  (
    .I0(SHADOW_CBE4),
    .I1(OUT_SEL64),
    .O(\PCI-CBE64/IO0/$1I2296/M1 )
  );
  X_OR2   \PCI-CBE64/IO0/$1I2296/$1I8  (
    .I0(\PCI-CBE64/IO0/$1I2296/M1 ),
    .I1(\PCI-CBE64/IO0/$1I2296/M0 ),
    .O(\PCI-CBE64/IO0/D_SLO )
  );
  X_AND2   \PCI-CBE64/IO0/$1I2296/$1I7  (
    .I0(\NlwInverterSignal_PCI-CBE64/IO0/$1I2296/$1I7/I0 ),
    .I1(M_CBE_INT4),
    .O(\PCI-CBE64/IO0/$1I2296/M0 )
  );
  X_AND2   \PCI-CBE64/IO0/$1I2303/$1I9  (
    .I0(\PCI-CBE64/$1N2781 ),
    .I1(\PCI-CBE64/IO0/$1N2321 ),
    .O(\PCI-CBE64/IO0/$1I2303/M1 )
  );
  X_OR2   \PCI-CBE64/IO0/$1I2303/$1I8  (
    .I0(\PCI-CBE64/IO0/$1I2303/M1 ),
    .I1(\PCI-CBE64/IO0/$1I2303/M0 ),
    .O(CBEOUT4)
  );
  X_AND2   \PCI-CBE64/IO0/$1I2303/$1I7  (
    .I0(\NlwInverterSignal_PCI-CBE64/IO0/$1I2303/$1I7/I0 ),
    .I1(\PCI-CBE64/IO0/D_SLO ),
    .O(\PCI-CBE64/IO0/$1I2303/M0 )
  );
  X_ZERO   \PCI-CBE64/$1I2777/$1I2218  (
    .O(\PCI-CBE64/$1I2777/$1N2216 )
  );
  X_BUF   \PCI-CBE64/$1I2777/L  (
    .I(\PCI-CBE64/$1I2777/$1N2216 ),
    .O(\PCI-CBE64/$1N2779 )
  );
  X_ZERO   \PCI-CBE64/$1I2780/$1I2218  (
    .O(\PCI-CBE64/$1I2780/$1N2216 )
  );
  X_BUF   \PCI-CBE64/$1I2780/L  (
    .I(\PCI-CBE64/$1I2780/$1N2216 ),
    .O(\PCI-CBE64/$1N2781 )
  );
  X_ZERO   \PCI-CBE64/$1I2782/$1I2218  (
    .O(\PCI-CBE64/$1I2782/$1N2216 )
  );
  X_BUF   \PCI-CBE64/$1I2782/L  (
    .I(\PCI-CBE64/$1I2782/$1N2216 ),
    .O(\PCI-CBE64/$1N2783 )
  );
  X_ZERO   \PCI-CBE64/$1I2784/$1I2218  (
    .O(\PCI-CBE64/$1I2784/$1N2216 )
  );
  X_BUF   \PCI-CBE64/$1I2784/L  (
    .I(\PCI-CBE64/$1I2784/$1N2216 ),
    .O(\PCI-CBE64/$1N2785 )
  );
  X_ZERO   \PCI-CBE64/$1I2786/$1I2218  (
    .O(\PCI-CBE64/$1I2786/$1N2216 )
  );
  X_BUF   \PCI-CBE64/$1I2786/L  (
    .I(\PCI-CBE64/$1I2786/$1N2216 ),
    .O(\PCI-CBE64/$1N2787 )
  );
  X_ZERO   \PCI-CBE64/$1I2788/$1I2218  (
    .O(\PCI-CBE64/$1I2788/$1N2216 )
  );
  X_BUF   \PCI-CBE64/$1I2788/L  (
    .I(\PCI-CBE64/$1I2788/$1N2216 ),
    .O(\PCI-CBE64/$1N2789 )
  );
  X_ZERO   \PCI-CBE64/$1I2790/$1I2218  (
    .O(\PCI-CBE64/$1I2790/$1N2216 )
  );
  X_BUF   \PCI-CBE64/$1I2790/L  (
    .I(\PCI-CBE64/$1I2790/$1N2216 ),
    .O(\PCI-CBE64/$1N2791 )
  );
  X_ZERO   \PCI-CBE64/$1I2792/$1I2218  (
    .O(\PCI-CBE64/$1I2792/$1N2216 )
  );
  X_BUF   \PCI-CBE64/$1I2792/L  (
    .I(\PCI-CBE64/$1I2792/$1N2216 ),
    .O(\PCI-CBE64/$1N2793 )
  );
  X_ZERO   \PCI-CBE64/$1I2794/$1I2218  (
    .O(\PCI-CBE64/$1I2794/$1N2216 )
  );
  X_BUF   \PCI-CBE64/$1I2794/L  (
    .I(\PCI-CBE64/$1I2794/$1N2216 ),
    .O(\PCI-CBE64/$1N2795 )
  );
  X_ZERO   \PCI-CBE64/$1I2796/$1I2218  (
    .O(\PCI-CBE64/$1I2796/$1N2216 )
  );
  X_BUF   \PCI-CBE64/$1I2796/L  (
    .I(\PCI-CBE64/$1I2796/$1N2216 ),
    .O(\PCI-CBE64/$1N2797 )
  );
  X_ZERO   \PCI-CBE64/$1I2798/$1I2218  (
    .O(\PCI-CBE64/$1I2798/$1N2216 )
  );
  X_BUF   \PCI-CBE64/$1I2798/L  (
    .I(\PCI-CBE64/$1I2798/$1N2216 ),
    .O(\PCI-CBE64/$1N2799 )
  );
  X_ZERO   \PCI-CBE64/$1I2800/$1I2218  (
    .O(\PCI-CBE64/$1I2800/$1N2216 )
  );
  X_BUF   \PCI-CBE64/$1I2800/L  (
    .I(\PCI-CBE64/$1I2800/$1N2216 ),
    .O(\PCI-CBE64/$1N2801 )
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD64/UPPER/Q15  (
    .CE(SHADOW_CE64),
    .CLK(CLK),
    .I(ADIO63),
    .O(SHADOW63),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD64/UPPER/Q9  (
    .CE(SHADOW_CE64),
    .CLK(CLK),
    .I(ADIO57),
    .O(SHADOW57),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD64/UPPER/Q13  (
    .CE(SHADOW_CE64),
    .CLK(CLK),
    .I(ADIO61),
    .O(SHADOW61),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD64/UPPER/Q10  (
    .CE(SHADOW_CE64),
    .CLK(CLK),
    .I(ADIO58),
    .O(SHADOW58),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD64/UPPER/Q14  (
    .CE(SHADOW_CE64),
    .CLK(CLK),
    .I(ADIO62),
    .O(SHADOW62),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD64/UPPER/Q12  (
    .CE(SHADOW_CE64),
    .CLK(CLK),
    .I(ADIO60),
    .O(SHADOW60),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD64/UPPER/Q11  (
    .CE(SHADOW_CE64),
    .CLK(CLK),
    .I(ADIO59),
    .O(SHADOW59),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD64/UPPER/Q8  (
    .CE(SHADOW_CE64),
    .CLK(CLK),
    .I(ADIO56),
    .O(SHADOW56),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD64/UPPER/Q7  (
    .CE(SHADOW_CE64),
    .CLK(CLK),
    .I(ADIO55),
    .O(SHADOW55),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD64/UPPER/Q1  (
    .CE(SHADOW_CE64),
    .CLK(CLK),
    .I(ADIO49),
    .O(SHADOW49),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD64/UPPER/Q5  (
    .CE(SHADOW_CE64),
    .CLK(CLK),
    .I(ADIO53),
    .O(SHADOW53),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD64/UPPER/Q3  (
    .CE(SHADOW_CE64),
    .CLK(CLK),
    .I(ADIO51),
    .O(SHADOW51),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD64/UPPER/Q0  (
    .CE(SHADOW_CE64),
    .CLK(CLK),
    .I(ADIO48),
    .O(SHADOW48),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD64/UPPER/Q2  (
    .CE(SHADOW_CE64),
    .CLK(CLK),
    .I(ADIO50),
    .O(SHADOW50),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD64/UPPER/Q4  (
    .CE(SHADOW_CE64),
    .CLK(CLK),
    .I(ADIO52),
    .O(SHADOW52),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD64/UPPER/Q6  (
    .CE(SHADOW_CE64),
    .CLK(CLK),
    .I(ADIO54),
    .O(SHADOW54),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD64/LOWER/Q15  (
    .CE(SHADOW_CE64),
    .CLK(CLK),
    .I(ADIO47),
    .O(SHADOW47),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD64/LOWER/Q9  (
    .CE(SHADOW_CE64),
    .CLK(CLK),
    .I(ADIO41),
    .O(SHADOW41),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD64/LOWER/Q13  (
    .CE(SHADOW_CE64),
    .CLK(CLK),
    .I(ADIO45),
    .O(SHADOW45),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD64/LOWER/Q10  (
    .CE(SHADOW_CE64),
    .CLK(CLK),
    .I(ADIO42),
    .O(SHADOW42),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD64/LOWER/Q14  (
    .CE(SHADOW_CE64),
    .CLK(CLK),
    .I(ADIO46),
    .O(SHADOW46),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD64/LOWER/Q12  (
    .CE(SHADOW_CE64),
    .CLK(CLK),
    .I(ADIO44),
    .O(SHADOW44),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD64/LOWER/Q11  (
    .CE(SHADOW_CE64),
    .CLK(CLK),
    .I(ADIO43),
    .O(SHADOW43),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD64/LOWER/Q8  (
    .CE(SHADOW_CE64),
    .CLK(CLK),
    .I(ADIO40),
    .O(SHADOW40),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD64/LOWER/Q7  (
    .CE(SHADOW_CE64),
    .CLK(CLK),
    .I(ADIO39),
    .O(SHADOW39),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD64/LOWER/Q1  (
    .CE(SHADOW_CE64),
    .CLK(CLK),
    .I(ADIO33),
    .O(SHADOW33),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD64/LOWER/Q5  (
    .CE(SHADOW_CE64),
    .CLK(CLK),
    .I(ADIO37),
    .O(SHADOW37),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD64/LOWER/Q3  (
    .CE(SHADOW_CE64),
    .CLK(CLK),
    .I(ADIO35),
    .O(SHADOW35),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD64/LOWER/Q0  (
    .CE(SHADOW_CE64),
    .CLK(CLK),
    .I(ADIO32),
    .O(SHADOW32),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD64/LOWER/Q2  (
    .CE(SHADOW_CE64),
    .CLK(CLK),
    .I(ADIO34),
    .O(SHADOW34),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD64/LOWER/Q4  (
    .CE(SHADOW_CE64),
    .CLK(CLK),
    .I(ADIO36),
    .O(SHADOW36),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD64/LOWER/Q6  (
    .CE(SHADOW_CE64),
    .CLK(CLK),
    .I(ADIO38),
    .O(SHADOW38),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD_CBE64/Q1  (
    .CE(SHADOW_CE64),
    .CLK(CLK),
    .I(M_CBE_INT5),
    .O(SHADOW_CBE5),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD_CBE64/Q3  (
    .CE(SHADOW_CE64),
    .CLK(CLK),
    .I(M_CBE_INT7),
    .O(SHADOW_CBE7),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD_CBE64/Q0  (
    .CE(SHADOW_CE64),
    .CLK(CLK),
    .I(M_CBE_INT4),
    .O(SHADOW_CBE4),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \SHD_CBE64/Q2  (
    .CE(SHADOW_CE64),
    .CLK(CLK),
    .I(M_CBE_INT6),
    .O(SHADOW_CBE6),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \FAIL_ADH/UPPER/Q15  (
    .CE(M_FIRST),
    .CLK(CLK),
    .I(ADIO63),
    .O(FAIL_ADH63),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \FAIL_ADH/UPPER/Q9  (
    .CE(M_FIRST),
    .CLK(CLK),
    .I(ADIO57),
    .O(FAIL_ADH57),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \FAIL_ADH/UPPER/Q13  (
    .CE(M_FIRST),
    .CLK(CLK),
    .I(ADIO61),
    .O(FAIL_ADH61),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \FAIL_ADH/UPPER/Q10  (
    .CE(M_FIRST),
    .CLK(CLK),
    .I(ADIO58),
    .O(FAIL_ADH58),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \FAIL_ADH/UPPER/Q14  (
    .CE(M_FIRST),
    .CLK(CLK),
    .I(ADIO62),
    .O(FAIL_ADH62),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \FAIL_ADH/UPPER/Q12  (
    .CE(M_FIRST),
    .CLK(CLK),
    .I(ADIO60),
    .O(FAIL_ADH60),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \FAIL_ADH/UPPER/Q11  (
    .CE(M_FIRST),
    .CLK(CLK),
    .I(ADIO59),
    .O(FAIL_ADH59),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \FAIL_ADH/UPPER/Q8  (
    .CE(M_FIRST),
    .CLK(CLK),
    .I(ADIO56),
    .O(FAIL_ADH56),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \FAIL_ADH/UPPER/Q7  (
    .CE(M_FIRST),
    .CLK(CLK),
    .I(ADIO55),
    .O(FAIL_ADH55),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \FAIL_ADH/UPPER/Q1  (
    .CE(M_FIRST),
    .CLK(CLK),
    .I(ADIO49),
    .O(FAIL_ADH49),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \FAIL_ADH/UPPER/Q5  (
    .CE(M_FIRST),
    .CLK(CLK),
    .I(ADIO53),
    .O(FAIL_ADH53),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \FAIL_ADH/UPPER/Q3  (
    .CE(M_FIRST),
    .CLK(CLK),
    .I(ADIO51),
    .O(FAIL_ADH51),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \FAIL_ADH/UPPER/Q0  (
    .CE(M_FIRST),
    .CLK(CLK),
    .I(ADIO48),
    .O(FAIL_ADH48),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \FAIL_ADH/UPPER/Q2  (
    .CE(M_FIRST),
    .CLK(CLK),
    .I(ADIO50),
    .O(FAIL_ADH50),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \FAIL_ADH/UPPER/Q4  (
    .CE(M_FIRST),
    .CLK(CLK),
    .I(ADIO52),
    .O(FAIL_ADH52),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \FAIL_ADH/UPPER/Q6  (
    .CE(M_FIRST),
    .CLK(CLK),
    .I(ADIO54),
    .O(FAIL_ADH54),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \FAIL_ADH/LOWER/Q15  (
    .CE(M_FIRST),
    .CLK(CLK),
    .I(ADIO47),
    .O(FAIL_ADH47),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \FAIL_ADH/LOWER/Q9  (
    .CE(M_FIRST),
    .CLK(CLK),
    .I(ADIO41),
    .O(FAIL_ADH41),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \FAIL_ADH/LOWER/Q13  (
    .CE(M_FIRST),
    .CLK(CLK),
    .I(ADIO45),
    .O(FAIL_ADH45),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \FAIL_ADH/LOWER/Q10  (
    .CE(M_FIRST),
    .CLK(CLK),
    .I(ADIO42),
    .O(FAIL_ADH42),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \FAIL_ADH/LOWER/Q14  (
    .CE(M_FIRST),
    .CLK(CLK),
    .I(ADIO46),
    .O(FAIL_ADH46),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \FAIL_ADH/LOWER/Q12  (
    .CE(M_FIRST),
    .CLK(CLK),
    .I(ADIO44),
    .O(FAIL_ADH44),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \FAIL_ADH/LOWER/Q11  (
    .CE(M_FIRST),
    .CLK(CLK),
    .I(ADIO43),
    .O(FAIL_ADH43),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \FAIL_ADH/LOWER/Q8  (
    .CE(M_FIRST),
    .CLK(CLK),
    .I(ADIO40),
    .O(FAIL_ADH40),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \FAIL_ADH/LOWER/Q7  (
    .CE(M_FIRST),
    .CLK(CLK),
    .I(ADIO39),
    .O(FAIL_ADH39),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \FAIL_ADH/LOWER/Q1  (
    .CE(M_FIRST),
    .CLK(CLK),
    .I(ADIO33),
    .O(FAIL_ADH33),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \FAIL_ADH/LOWER/Q5  (
    .CE(M_FIRST),
    .CLK(CLK),
    .I(ADIO37),
    .O(FAIL_ADH37),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \FAIL_ADH/LOWER/Q3  (
    .CE(M_FIRST),
    .CLK(CLK),
    .I(ADIO35),
    .O(FAIL_ADH35),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \FAIL_ADH/LOWER/Q0  (
    .CE(M_FIRST),
    .CLK(CLK),
    .I(ADIO32),
    .O(FAIL_ADH32),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \FAIL_ADH/LOWER/Q2  (
    .CE(M_FIRST),
    .CLK(CLK),
    .I(ADIO34),
    .O(FAIL_ADH34),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \FAIL_ADH/LOWER/Q4  (
    .CE(M_FIRST),
    .CLK(CLK),
    .I(ADIO36),
    .O(FAIL_ADH36),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \FAIL_ADH/LOWER/Q6  (
    .CE(M_FIRST),
    .CLK(CLK),
    .I(ADIO38),
    .O(FAIL_ADH38),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \FAIL_CBH/Q1  (
    .CE(M_FIRST),
    .CLK(CLK),
    .I(M_CBE_INT5),
    .O(FAIL_CBH5),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \FAIL_CBH/Q3  (
    .CE(M_FIRST),
    .CLK(CLK),
    .I(M_CBE_INT7),
    .O(FAIL_CBH7),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \FAIL_CBH/Q0  (
    .CE(M_FIRST),
    .CLK(CLK),
    .I(M_CBE_INT4),
    .O(FAIL_CBH4),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_FF #(
    .INIT ( 1'b0 ))
  \FAIL_CBH/Q2  (
    .CE(M_FIRST),
    .CLK(CLK),
    .I(M_CBE_INT6),
    .O(FAIL_CBH6),
    .RST(NlwRenamedSig_OI_RST),
    .SET(GND)
  );
  X_INV   \NlwInverterBlock_$3I3487/I0  (
    .I(CFG0),
    .O(\NlwInverterSignal_$3I3487/I0 )
  );
  X_INV   \NlwInverterBlock_$3I3492/I0  (
    .I(CFG37),
    .O(\NlwInverterSignal_$3I3492/I0 )
  );
  X_INV   \NlwInverterBlock_$3I3496/I0  (
    .I(CFG74),
    .O(\NlwInverterSignal_$3I3496/I0 )
  );
  X_INV   \NlwInverterBlock_$4I4017/I0  (
    .I(INTR_N),
    .O(\NlwInverterSignal_$4I4017/I0 )
  );
  X_INV   \NlwInverterBlock_$4I4017/I1  (
    .I(NlwRenamedSig_OI_CSR10),
    .O(\NlwInverterSignal_$4I4017/I1 )
  );
  X_INV   \NlwInverterBlock_$4I4017/O  (
    .I(\NlwInverterSignal_$4I4017/O ),
    .O(OE_INTA)
  );
  X_INV   \NlwInverterBlock_$6I1168/I0  (
    .I(CFG240),
    .O(\NlwInverterSignal_$6I1168/I0 )
  );
  X_INV   \NlwInverterBlock_$6I1168/I1  (
    .I(CFG110),
    .O(\NlwInverterSignal_$6I1168/I1 )
  );
  X_INV   \NlwInverterBlock_$6I1169/I0  (
    .I(CFG73),
    .O(\NlwInverterSignal_$6I1169/I0 )
  );
  X_INV   \NlwInverterBlock_$6I1170/I0  (
    .I(CFG240),
    .O(\NlwInverterSignal_$6I1170/I0 )
  );
  X_INV   \NlwInverterBlock_$6I1172/I0  (
    .I(CFG36),
    .O(\NlwInverterSignal_$6I1172/I0 )
  );
  X_INV   \NlwInverterBlock_$7I129/I0  (
    .I(\TRDY- ),
    .O(\NlwInverterSignal_$7I129/I0 )
  );
  X_INV   \NlwInverterBlock_$7I129/I1  (
    .I(\IRDY- ),
    .O(\NlwInverterSignal_$7I129/I1 )
  );
  X_INV   \NlwInverterBlock_$7I130/I0  (
    .I(\TRDY- ),
    .O(\NlwInverterSignal_$7I130/I0 )
  );
  X_INV   \NlwInverterBlock_$7I131/I0  (
    .I(\STOP- ),
    .O(\NlwInverterSignal_$7I131/I0 )
  );
  X_INV   \NlwInverterBlock_$7I132/I0  (
    .I(\DEVSEL- ),
    .O(\NlwInverterSignal_$7I132/I0 )
  );
  X_INV   \NlwInverterBlock_$7I132/I1  (
    .I(\STOP- ),
    .O(\NlwInverterSignal_$7I132/I1 )
  );
  X_INV   \NlwInverterBlock_$7I133/I0  (
    .I(\DEVSEL- ),
    .O(\NlwInverterSignal_$7I133/I0 )
  );
  X_INV   \NlwInverterBlock_$7I133/I1  (
    .I(\STOP- ),
    .O(\NlwInverterSignal_$7I133/I1 )
  );
  X_INV   \NlwInverterBlock_$7I133/I2  (
    .I(\TRDY- ),
    .O(\NlwInverterSignal_$7I133/I2 )
  );
  X_INV   \NlwInverterBlock_$7I134/I0  (
    .I(\STOP- ),
    .O(\NlwInverterSignal_$7I134/I0 )
  );
  X_INV   \NlwInverterBlock_$7I141/I0  (
    .I(\STOP- ),
    .O(\NlwInverterSignal_$7I141/I0 )
  );
  X_INV   \NlwInverterBlock_$7I141/I1  (
    .I(\TRDY- ),
    .O(\NlwInverterSignal_$7I141/I1 )
  );
  X_ONE   NlwBlock_PCI_LC_I_VCC (
    .O(VCC)
  );
  X_ZERO   NlwBlock_PCI_LC_I_GND (
    .O(GND)
  );
  X_INV   \NlwInverterBlock_$7I863/I0  (
    .I(EX),
    .O(\NlwInverterSignal_$7I863/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/$4I3271/I0  (
    .I(NlwRenamedSig_OI_OE_CBE64),
    .O(\NlwInverterSignal_MASTER/$4I3271/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/$4I3271/I1  (
    .I(M_WRDN),
    .O(\NlwInverterSignal_MASTER/$4I3271/I1 )
  );
  X_INV   \NlwInverterBlock_MASTER/$4I3271/I2  (
    .I(\IIRDY_I- ),
    .O(\NlwInverterSignal_MASTER/$4I3271/I2 )
  );
  X_INV   \NlwInverterBlock_MASTER/$4I3102/I0  (
    .I(FAIL64_INT),
    .O(\NlwInverterSignal_MASTER/$4I3102/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/$4I3102/I1  (
    .I(\TRDY- ),
    .O(\NlwInverterSignal_MASTER/$4I3102/I1 )
  );
  X_INV   \NlwInverterBlock_MASTER/$4I3072/I0  (
    .I(\MASTER/$4N3030 ),
    .O(\NlwInverterSignal_MASTER/$4I3072/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/$4I3051/I0  (
    .I(\STOP- ),
    .O(\NlwInverterSignal_MASTER/$4I3051/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/$4I2686/I0  (
    .I(\MASTER/IIRDY- ),
    .O(\NlwInverterSignal_MASTER/$4I2686/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/$4I2686/I1  (
    .I(\TRDY- ),
    .O(\NlwInverterSignal_MASTER/$4I2686/I1 )
  );
  X_INV   \NlwInverterBlock_MASTER/$4I2686/I2  (
    .I(M_WRDN),
    .O(\NlwInverterSignal_MASTER/$4I2686/I2 )
  );
  X_INV   \NlwInverterBlock_MASTER/I_IDLE/$1I2807/I0  (
    .I(ADDR_BE),
    .O(\NlwInverterSignal_MASTER/I_IDLE/$1I2807/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/I_IDLE/$1I2715/I0  (
    .I(GNT_IN),
    .O(\NlwInverterSignal_MASTER/I_IDLE/$1I2715/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/I_IDLE/$1I2715/I1  (
    .I(\GNT- ),
    .O(\NlwInverterSignal_MASTER/I_IDLE/$1I2715/I1 )
  );
  X_INV   \NlwInverterBlock_MASTER/I_IDLE/$1I2715/O  (
    .I(\NlwInverterSignal_MASTER/I_IDLE/$1I2715/O ),
    .O(\MASTER/I_IDLE/ADDR_GNT )
  );
  X_INV   \NlwInverterBlock_MASTER/I_IDLE/$1I2647/I0  (
    .I(\MASTER/IFRAME- ),
    .O(\NlwInverterSignal_MASTER/I_IDLE/$1I2647/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/I_IDLE/$1I2594/I0  (
    .I(\MASTER/DEV_TO ),
    .O(\NlwInverterSignal_MASTER/I_IDLE/$1I2594/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/I_IDLE/$1I2593/I0  (
    .I(\MASTER/I_IDLE/M_DATA_C2 ),
    .O(\NlwInverterSignal_MASTER/I_IDLE/$1I2593/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/ADDR/$1I2632/I0  (
    .I(GNT_IN),
    .O(\NlwInverterSignal_MASTER/ADDR/$1I2632/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/ADDR/$1I2630/O  (
    .I(\NlwInverterSignal_MASTER/ADDR/$1I2630/O ),
    .O(\MASTER/ADDR/NS_MAN )
  );
  X_INV   \NlwInverterBlock_MASTER/ADDR/$1I2623/I0  (
    .I(ADDR_BE),
    .O(\NlwInverterSignal_MASTER/ADDR/$1I2623/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/ADDR/$1I2602/I0  (
    .I(GNT_IN),
    .O(\NlwInverterSignal_MASTER/ADDR/$1I2602/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/DR_BUS/$1I2913/I0  (
    .I(\MASTER/DR_BUS/BBBRGH ),
    .O(\NlwInverterSignal_MASTER/DR_BUS/$1I2913/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/DR_BUS/$1I2913/I1  (
    .I(\GNT- ),
    .O(\NlwInverterSignal_MASTER/DR_BUS/$1I2913/I1 )
  );
  X_INV   \NlwInverterBlock_MASTER/DR_BUS/$1I2913/I2  (
    .I(ADDR_BE),
    .O(\NlwInverterSignal_MASTER/DR_BUS/$1I2913/I2 )
  );
  X_INV   \NlwInverterBlock_MASTER/DR_BUS/$1I2805/I0  (
    .I(\MASTER/M_ENABLE ),
    .O(\NlwInverterSignal_MASTER/DR_BUS/$1I2805/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/DR_BUS/$1I2805/I1  (
    .I(\MASTER/REQUEST ),
    .O(\NlwInverterSignal_MASTER/DR_BUS/$1I2805/I1 )
  );
  X_INV   \NlwInverterBlock_MASTER/DR_BUS/$1I2787/I0  (
    .I(\GNT- ),
    .O(\NlwInverterSignal_MASTER/DR_BUS/$1I2787/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/DR_BUS/$1I2752/I0  (
    .I(\GNT- ),
    .O(\NlwInverterSignal_MASTER/DR_BUS/$1I2752/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/DR_BUS/$1I2752/I1  (
    .I(\MASTER/REQUEST ),
    .O(\NlwInverterSignal_MASTER/DR_BUS/$1I2752/I1 )
  );
  X_INV   \NlwInverterBlock_MASTER/DR_BUS/$1I2732/I0  (
    .I(ADDR_BE),
    .O(\NlwInverterSignal_MASTER/DR_BUS/$1I2732/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/DR_BUS/$1I2732/I1  (
    .I(\GNT- ),
    .O(\NlwInverterSignal_MASTER/DR_BUS/$1I2732/I1 )
  );
  X_INV   \NlwInverterBlock_MASTER/DR_BUS/$1I2721/I0  (
    .I(\MASTER/DR_BUS/COND ),
    .O(\NlwInverterSignal_MASTER/DR_BUS/$1I2721/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/DR_BUS/$1I2719/I0  (
    .I(\MASTER/IFRAME- ),
    .O(\NlwInverterSignal_MASTER/DR_BUS/$1I2719/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/DR_BUS/$1I2706/I0  (
    .I(\MASTER/DEV_TO ),
    .O(\NlwInverterSignal_MASTER/DR_BUS/$1I2706/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/DR_BUS/$1I2704/I0  (
    .I(\GNT- ),
    .O(\NlwInverterSignal_MASTER/DR_BUS/$1I2704/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/DR_BUS/$1I2908/$1I7/I0  (
    .I(\$1N4834 ),
    .O(\NlwInverterSignal_MASTER/DR_BUS/$1I2908/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/DR_BUS/$1I2917/$1I7/I0  (
    .I(\$1N4834 ),
    .O(\NlwInverterSignal_MASTER/DR_BUS/$1I2917/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/M_DATA/$1I2590/I0  (
    .I(GNT_IN),
    .O(\NlwInverterSignal_MASTER/M_DATA/$1I2590/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/M_DATA/$1I2518/I0  (
    .I(\MASTER/IFRAME- ),
    .O(\NlwInverterSignal_MASTER/M_DATA/$1I2518/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/M_DATA/$1I2502/I0  (
    .I(\MASTER/DEV_TO ),
    .O(\NlwInverterSignal_MASTER/M_DATA/$1I2502/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/$1I2914/$1I2947/I0  (
    .I(\MASTER/M_ENABLE ),
    .O(\NlwInverterSignal_MASTER/$1I2914/$1I2947/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/$1I2914/$1I2931/I0  (
    .I(\MASTER/$1I2914/LOCKOUT ),
    .O(\NlwInverterSignal_MASTER/$1I2914/$1I2931/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/$1I2914/$1I2927/I0  (
    .I(M_DATA_INT),
    .O(\NlwInverterSignal_MASTER/$1I2914/$1I2927/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/$1I2914/$1I2908/I0  (
    .I(M_DATA_INT),
    .O(\NlwInverterSignal_MASTER/$1I2914/$1I2908/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/$1I2914/$1I2895/I0  (
    .I(\MASTER/$1I2914/LOCKOUT ),
    .O(\NlwInverterSignal_MASTER/$1I2914/$1I2895/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/$1I2914/$1I2880/I0  (
    .I(M_DATA_INT),
    .O(\NlwInverterSignal_MASTER/$1I2914/$1I2880/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/$1I2914/$1I2879/I0  (
    .I(\MASTER/$1I2914/LOCKOUT ),
    .O(\NlwInverterSignal_MASTER/$1I2914/$1I2879/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/$1I2914/$1I2853/$1I2213/I0  (
    .I(\MASTER/$1I2914/CANCEL ),
    .O(\NlwInverterSignal_MASTER/$1I2914/$1I2853/$1I2213/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/$1I2914/$1I2864/$1I2213/I0  (
    .I(\MASTER/$1I2914/CANCEL ),
    .O(\NlwInverterSignal_MASTER/$1I2914/$1I2864/$1I2213/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/$1I2914/$1I2932/$1I2213/I0  (
    .I(\MASTER/$1I2914/END_OF_XFER ),
    .O(\NlwInverterSignal_MASTER/$1I2914/$1I2932/$1I2213/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/FRAME/$2I3528/I0  (
    .I(\STOP- ),
    .O(\NlwInverterSignal_MASTER/FRAME/$2I3528/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/FRAME/$2I3511/I0  (
    .I(\STOP- ),
    .O(\NlwInverterSignal_MASTER/FRAME/$2I3511/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/FRAME/$2I3464/I0  (
    .I(\MASTER/FRAME/$2N3475 ),
    .O(\NlwInverterSignal_MASTER/FRAME/$2I3464/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/FRAME/$2I3463/I0  (
    .I(\MASTER/FRAME/$2N3449 ),
    .O(\NlwInverterSignal_MASTER/FRAME/$2I3463/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/FRAME/$1I3470/O  (
    .I(\NlwInverterSignal_MASTER/FRAME/$1I3470/O ),
    .O(\MASTER/FRAME/NS_S_1 )
  );
  X_INV   \NlwInverterBlock_MASTER/FRAME/$1I3466/I0  (
    .I(GNT_IN),
    .O(\NlwInverterSignal_MASTER/FRAME/$1I3466/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/FRAME/$1I3393/I0  (
    .I(M_READY),
    .O(\NlwInverterSignal_MASTER/FRAME/$1I3393/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/FRAME/$1I3368/O  (
    .I(\NlwInverterSignal_MASTER/FRAME/$1I3368/O ),
    .O(\MASTER/FRAME/NS_S_0 )
  );
  X_INV   \NlwInverterBlock_MASTER/FRAME/$1I3323/I0  (
    .I(TRDY_M),
    .O(\NlwInverterSignal_MASTER/FRAME/$1I3323/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/FRAME/$1I3323/O  (
    .I(\NlwInverterSignal_MASTER/FRAME/$1I3323/O ),
    .O(FRAME_CE)
  );
  X_INV   \NlwInverterBlock_MASTER/FRAME/$1I3322/I0  (
    .I(\IIRDY_I- ),
    .O(\NlwInverterSignal_MASTER/FRAME/$1I3322/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/FRAME/$1I3144/I0  (
    .I(\MASTER/DEV_TO ),
    .O(\NlwInverterSignal_MASTER/FRAME/$1I3144/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/FRAME/$1I3144/I1  (
    .I(\IFRAME_I- ),
    .O(\NlwInverterSignal_MASTER/FRAME/$1I3144/I1 )
  );
  X_INV   \NlwInverterBlock_MASTER/FRAME/$1I3144/I2  (
    .I(FAIL64_INT),
    .O(\NlwInverterSignal_MASTER/FRAME/$1I3144/I2 )
  );
  X_INV   \NlwInverterBlock_MASTER/FRAME/$1I3467/$1I7/I0  (
    .I(TRDY_M),
    .O(\NlwInverterSignal_MASTER/FRAME/$1I3467/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/FRAME/$2I3559/$1I7/I0  (
    .I(CFG254),
    .O(\NlwInverterSignal_MASTER/FRAME/$2I3559/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/IRDY/$2I3437/I0  (
    .I(\IFRAME_I- ),
    .O(\NlwInverterSignal_MASTER/IRDY/$2I3437/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/IRDY/$2I3435/O  (
    .I(\NlwInverterSignal_MASTER/IRDY/$2I3435/O ),
    .O(\MASTER/IRDY/$2N3355 )
  );
  X_INV   \NlwInverterBlock_MASTER/IRDY/$2I3390/O  (
    .I(\NlwInverterSignal_MASTER/IRDY/$2I3390/O ),
    .O(\MASTER/IRDY/$2N3385 )
  );
  X_INV   \NlwInverterBlock_MASTER/IRDY/$2I3332/I0  (
    .I(TRDY_M),
    .O(\NlwInverterSignal_MASTER/IRDY/$2I3332/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/IRDY/$2I3332/O  (
    .I(\NlwInverterSignal_MASTER/IRDY/$2I3332/O ),
    .O(\MASTER/IRDY/$2N3294 )
  );
  X_INV   \NlwInverterBlock_MASTER/IRDY/$2I3233/I0  (
    .I(M_DATA_INT),
    .O(\NlwInverterSignal_MASTER/IRDY/$2I3233/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/IRDY/$1I3779/I0  (
    .I(\IFRAME_I- ),
    .O(\NlwInverterSignal_MASTER/IRDY/$1I3779/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/IRDY/$1I3779/O  (
    .I(\NlwInverterSignal_MASTER/IRDY/$1I3779/O ),
    .O(\MASTER/IRDY/NS_0 )
  );
  X_INV   \NlwInverterBlock_MASTER/IRDY/$1I3738/I0  (
    .I(\IFRAME_I- ),
    .O(\NlwInverterSignal_MASTER/IRDY/$1I3738/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/IRDY/$1I3738/I1  (
    .I(\MASTER/DEV_TO ),
    .O(\NlwInverterSignal_MASTER/IRDY/$1I3738/I1 )
  );
  X_INV   \NlwInverterBlock_MASTER/IRDY/$1I3699/I0  (
    .I(\MASTER/IFRAME- ),
    .O(\NlwInverterSignal_MASTER/IRDY/$1I3699/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/IRDY/$1I3698/I0  (
    .I(\MASTER/DEV_TO ),
    .O(\NlwInverterSignal_MASTER/IRDY/$1I3698/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/IRDY/$1I3498/I0  (
    .I(\IIRDY_I- ),
    .O(\NlwInverterSignal_MASTER/IRDY/$1I3498/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/IRDY/$1I3491/I0  (
    .I(\IIRDY_I- ),
    .O(\NlwInverterSignal_MASTER/IRDY/$1I3491/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/IRDY/$1I3487/I0  (
    .I(TRDY_M),
    .O(\NlwInverterSignal_MASTER/IRDY/$1I3487/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/IRDY/$1I3487/O  (
    .I(\NlwInverterSignal_MASTER/IRDY/$1I3487/O ),
    .O(\MASTER/IRDY/CORE_READY )
  );
  X_INV   \NlwInverterBlock_MASTER/IRDY/$1I3211/O  (
    .I(\NlwInverterSignal_MASTER/IRDY/$1I3211/O ),
    .O(\MASTER/IRDY/NS_1 )
  );
  X_INV   \NlwInverterBlock_MASTER/IRDY/$1I3227/$1I7/I0  (
    .I(STOP_I),
    .O(\NlwInverterSignal_MASTER/IRDY/$1I3227/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/IRDY/$1I3492/$1I7/I0  (
    .I(ACK64_I),
    .O(\NlwInverterSignal_MASTER/IRDY/$1I3492/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/IRDY/$2I3285/$1I7/I0  (
    .I(STOP_I),
    .O(\NlwInverterSignal_MASTER/IRDY/$2I3285/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/REQ/$1I2726/O  (
    .I(\NlwInverterSignal_MASTER/REQ/$1I2726/O ),
    .O(\MASTER/REQ/S_TAR_OR )
  );
  X_INV   \NlwInverterBlock_MASTER/REQ/$1I2721/O  (
    .I(\NlwInverterSignal_MASTER/REQ/$1I2721/O ),
    .O(\MASTER/NS_REQ- )
  );
  X_INV   \NlwInverterBlock_MASTER/REQ/$1I2670/I0  (
    .I(\MASTER/REQ/M_DATA_Q ),
    .O(\NlwInverterSignal_MASTER/REQ/$1I2670/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/REQ/$1I2708/$1I2213/I0  (
    .I(\MASTER/REQ/SOXFER ),
    .O(\NlwInverterSignal_MASTER/REQ/$1I2708/$1I2213/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/REQ64/$2I3431/I0  (
    .I(\MASTER/REQ64/$2N3430 ),
    .O(\NlwInverterSignal_MASTER/REQ64/$2I3431/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/REQ64/$2I3411/I0  (
    .I(\STOP- ),
    .O(\NlwInverterSignal_MASTER/REQ64/$2I3411/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/REQ64/$2I3406/I0  (
    .I(\MASTER/REQ64/$2N3428 ),
    .O(\NlwInverterSignal_MASTER/REQ64/$2I3406/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/REQ64/$2I3393/I0  (
    .I(\STOP- ),
    .O(\NlwInverterSignal_MASTER/REQ64/$2I3393/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/REQ64/$1I3616/I0  (
    .I(GNT_IN),
    .O(\NlwInverterSignal_MASTER/REQ64/$1I3616/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/REQ64/$1I3614/I0  (
    .I(M_READY),
    .O(\NlwInverterSignal_MASTER/REQ64/$1I3614/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/REQ64/$1I3607/I0  (
    .I(\MASTER/DEV_TO ),
    .O(\NlwInverterSignal_MASTER/REQ64/$1I3607/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/REQ64/$1I3607/I1  (
    .I(\IREQ64_I- ),
    .O(\NlwInverterSignal_MASTER/REQ64/$1I3607/I1 )
  );
  X_INV   \NlwInverterBlock_MASTER/REQ64/$1I3607/I2  (
    .I(FAIL64_INT),
    .O(\NlwInverterSignal_MASTER/REQ64/$1I3607/I2 )
  );
  X_INV   \NlwInverterBlock_MASTER/REQ64/$1I3569/O  (
    .I(\NlwInverterSignal_MASTER/REQ64/$1I3569/O ),
    .O(\MASTER/REQ64/NS_S_0 )
  );
  X_INV   \NlwInverterBlock_MASTER/REQ64/$1I3561/O  (
    .I(\NlwInverterSignal_MASTER/REQ64/$1I3561/O ),
    .O(\MASTER/REQ64/NS_S_1 )
  );
  X_INV   \NlwInverterBlock_MASTER/REQ64/$1I3540/I0  (
    .I(\IIRDY_I- ),
    .O(\NlwInverterSignal_MASTER/REQ64/$1I3540/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/REQ64/$1I3534/I0  (
    .I(TRDY_M),
    .O(\NlwInverterSignal_MASTER/REQ64/$1I3534/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/REQ64/$1I3534/O  (
    .I(\NlwInverterSignal_MASTER/REQ64/$1I3534/O ),
    .O(REQ64_CE)
  );
  X_INV   \NlwInverterBlock_MASTER/REQ64/$1I3562/$1I7/I0  (
    .I(TRDY_M),
    .O(\NlwInverterSignal_MASTER/REQ64/$1I3562/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/REQ64/$2I3446/$1I7/I0  (
    .I(CFG254),
    .O(\NlwInverterSignal_MASTER/REQ64/$2I3446/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/XFERFAIL/$1I3024/I0  (
    .I(\IIRDY_I- ),
    .O(\NlwInverterSignal_MASTER/XFERFAIL/$1I3024/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/XFERFAIL/$1I3019/I0  (
    .I(DEVSEL_I),
    .O(\NlwInverterSignal_MASTER/XFERFAIL/$1I3019/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$8I4093/I0  (
    .I(\MASTER/OE_FRAME/OE_REQ64_INT_525 ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$8I4093/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$8I4047/O  (
    .I(\NlwInverterSignal_MASTER/OE_FRAME/$8I4047/O ),
    .O(\MASTER/OE_FRAME/NS_OER_0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$8I4045/I0  (
    .I(STOP_I),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$8I4045/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$8I4045/I1  (
    .I(TRDY_M),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$8I4045/I1 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$8I4044/I0  (
    .I(STOP_I),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$8I4044/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$8I4044/I1  (
    .I(TRDY_M),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$8I4044/I1 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$8I4043/O  (
    .I(\NlwInverterSignal_MASTER/OE_FRAME/$8I4043/O ),
    .O(\MASTER/OE_FRAME/$8N4018 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$8I4007/I0  (
    .I(\MASTER/OE_FRAME/OE_FRAME_INT_509 ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$8I4007/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$8I3975/O  (
    .I(\NlwInverterSignal_MASTER/OE_FRAME/$8I3975/O ),
    .O(\MASTER/OE_FRAME/$8N3992 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$8I3974/I0  (
    .I(STOP_I),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$8I3974/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$8I3974/I1  (
    .I(TRDY_M),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$8I3974/I1 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$8I3973/I0  (
    .I(STOP_I),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$8I3973/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$8I3973/I1  (
    .I(TRDY_M),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$8I3973/I1 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$8I3971/O  (
    .I(\NlwInverterSignal_MASTER/OE_FRAME/$8I3971/O ),
    .O(\MASTER/OE_FRAME/NS_OEF_0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$7I3977/O  (
    .I(\NlwInverterSignal_MASTER/OE_FRAME/$7I3977/O ),
    .O(\MASTER/OE_FRAME/NS64_1 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$7I3976/O  (
    .I(\NlwInverterSignal_MASTER/OE_FRAME/$7I3976/O ),
    .O(\MASTER/OE_FRAME/MISC64_2 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$7I3975/I0  (
    .I(GNT_IN),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$7I3975/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$7I3975/I1  (
    .I(\MASTER/OE_FRAME/DR_BUS1 ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$7I3975/I1 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$7I3968/I0  (
    .I(STOP_I),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$7I3968/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$7I3968/I1  (
    .I(TRDY_M),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$7I3968/I1 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$7I3966/I0  (
    .I(STOP_I),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$7I3966/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$7I3966/I1  (
    .I(TRDY_M),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$7I3966/I1 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$7I3965/O  (
    .I(\NlwInverterSignal_MASTER/OE_FRAME/$7I3965/O ),
    .O(\MASTER/OE_FRAME/$7N3936 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$6I3740/O  (
    .I(\NlwInverterSignal_MASTER/OE_FRAME/$6I3740/O ),
    .O(\MASTER/OE_FRAME/NS_1 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$6I3739/O  (
    .I(\NlwInverterSignal_MASTER/OE_FRAME/$6I3739/O ),
    .O(\MASTER/OE_FRAME/MISC_2 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$6I3738/I0  (
    .I(GNT_IN),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$6I3738/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$6I3738/I1  (
    .I(\MASTER/OE_FRAME/DR_BUS1 ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$6I3738/I1 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$6I3731/I0  (
    .I(STOP_I),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$6I3731/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$6I3731/I1  (
    .I(TRDY_M),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$6I3731/I1 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$6I3729/I0  (
    .I(STOP_I),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$6I3729/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$6I3729/I1  (
    .I(TRDY_M),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$6I3729/I1 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$6I3728/O  (
    .I(\NlwInverterSignal_MASTER/OE_FRAME/$6I3728/O ),
    .O(\MASTER/OE_FRAME/$6N3707 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$5I3899/I0  (
    .I(OE_AD_T_B64),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$5I3899/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$5I3899/O  (
    .I(\NlwInverterSignal_MASTER/OE_FRAME/$5I3899/O ),
    .O(\MASTER/OE_FRAME/$5N3897 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$5I3898/I0  (
    .I(\MASTER/OE_FRAME/$5N3897 ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$5I3898/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$5I3898/I1  (
    .I(EOT),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$5I3898/I1 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$5I3898/O  (
    .I(\NlwInverterSignal_MASTER/OE_FRAME/$5I3898/O ),
    .O(\MASTER/OE_FRAME/AD_B64 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$5I3893/I0  (
    .I(\MASTER/OE_FRAME/AD_T64 ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$5I3893/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$5I3893/O  (
    .I(\NlwInverterSignal_MASTER/OE_FRAME/$5I3893/O ),
    .O(\MASTER/OE_FRAME/$5N3892 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$5I3891/I0  (
    .I(EOT),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$5I3891/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$5I3891/O  (
    .I(\NlwInverterSignal_MASTER/OE_FRAME/$5I3891/O ),
    .O(\MASTER/OE_FRAME/CB64 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$5I3890/I0  (
    .I(\MASTER/OE_FRAME/CB64 ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$5I3890/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$5I3890/O  (
    .I(\NlwInverterSignal_MASTER/OE_FRAME/$5I3890/O ),
    .O(\MASTER/OE_FRAME/$5N3876 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$5I3889/I0  (
    .I(\MASTER/OE_FRAME/AD_LT64 ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$5I3889/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$5I3889/O  (
    .I(\NlwInverterSignal_MASTER/OE_FRAME/$5I3889/O ),
    .O(\MASTER/OE_FRAME/$5N3873 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$5I3888/I0  (
    .I(\MASTER/OE_FRAME/AD_LB64 ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$5I3888/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$5I3888/O  (
    .I(\NlwInverterSignal_MASTER/OE_FRAME/$5I3888/O ),
    .O(\MASTER/OE_FRAME/$5N3872 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$5I3887/I0  (
    .I(\MASTER/OE_FRAME/AD_B64 ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$5I3887/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$5I3887/O  (
    .I(\NlwInverterSignal_MASTER/OE_FRAME/$5I3887/O ),
    .O(\MASTER/OE_FRAME/$5N3871 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$5I3886/I0  (
    .I(OE_AD_T_LB64),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$5I3886/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$5I3886/O  (
    .I(\NlwInverterSignal_MASTER/OE_FRAME/$5I3886/O ),
    .O(\MASTER/OE_FRAME/$5N3896 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$5I3885/I0  (
    .I(OE_AD_T_LT64),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$5I3885/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$5I3885/O  (
    .I(\NlwInverterSignal_MASTER/OE_FRAME/$5I3885/O ),
    .O(\MASTER/OE_FRAME/$5N3895 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$5I3884/I0  (
    .I(OE_AD_T_T64),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$5I3884/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$5I3884/O  (
    .I(\NlwInverterSignal_MASTER/OE_FRAME/$5I3884/O ),
    .O(\MASTER/OE_FRAME/$5N3894 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$5I3883/I0  (
    .I(\MASTER/OE_FRAME/$5N3896 ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$5I3883/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$5I3883/I1  (
    .I(EOT),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$5I3883/I1 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$5I3883/O  (
    .I(\NlwInverterSignal_MASTER/OE_FRAME/$5I3883/O ),
    .O(\MASTER/OE_FRAME/AD_LB64 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$5I3882/I0  (
    .I(\MASTER/OE_FRAME/$5N3895 ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$5I3882/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$5I3882/I1  (
    .I(EOT),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$5I3882/I1 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$5I3882/O  (
    .I(\NlwInverterSignal_MASTER/OE_FRAME/$5I3882/O ),
    .O(\MASTER/OE_FRAME/AD_LT64 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$5I3881/I0  (
    .I(\MASTER/OE_FRAME/$5N3894 ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$5I3881/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$5I3881/I1  (
    .I(EOT),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$5I3881/I1 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$5I3881/O  (
    .I(\NlwInverterSignal_MASTER/OE_FRAME/$5I3881/O ),
    .O(\MASTER/OE_FRAME/AD_T64 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$4I3785/I0  (
    .I(EOT),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$4I3785/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$4I3785/O  (
    .I(\NlwInverterSignal_MASTER/OE_FRAME/$4I3785/O ),
    .O(\MASTER/OE_FRAME/CB32 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$4I3784/I0  (
    .I(\MASTER/OE_FRAME/CB32 ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$4I3784/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$4I3784/O  (
    .I(\NlwInverterSignal_MASTER/OE_FRAME/$4I3784/O ),
    .O(NlwRenamedSig_OI_OE_CBE)
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$4I3783/I0  (
    .I(\MASTER/OE_FRAME/AD_T ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$4I3783/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$4I3783/O  (
    .I(\NlwInverterSignal_MASTER/OE_FRAME/$4I3783/O ),
    .O(NlwRenamedSig_OI_OE_ADO_T)
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$4I3782/I0  (
    .I(\MASTER/OE_FRAME/AD_LT ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$4I3782/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$4I3782/O  (
    .I(\NlwInverterSignal_MASTER/OE_FRAME/$4I3782/O ),
    .O(NlwRenamedSig_OI_OE_ADO_LT)
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$4I3781/I0  (
    .I(\MASTER/OE_FRAME/AD_LB ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$4I3781/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$4I3781/O  (
    .I(\NlwInverterSignal_MASTER/OE_FRAME/$4I3781/O ),
    .O(NlwRenamedSig_OI_OE_ADO_LB)
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$4I3780/I0  (
    .I(\MASTER/OE_FRAME/AD_B ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$4I3780/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$4I3780/O  (
    .I(\NlwInverterSignal_MASTER/OE_FRAME/$4I3780/O ),
    .O(NlwRenamedSig_OI_OE_ADO_B)
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$4I3779/I0  (
    .I(\MASTER/OE_FRAME/$4N3741 ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$4I3779/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$4I3779/I1  (
    .I(EOT),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$4I3779/I1 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$4I3779/O  (
    .I(\NlwInverterSignal_MASTER/OE_FRAME/$4I3779/O ),
    .O(\MASTER/OE_FRAME/AD_B )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$4I3778/I0  (
    .I(OE_AD_T_B),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$4I3778/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$4I3778/O  (
    .I(\NlwInverterSignal_MASTER/OE_FRAME/$4I3778/O ),
    .O(\MASTER/OE_FRAME/$4N3741 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$4I3776/I0  (
    .I(OE_AD_T_LB),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$4I3776/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$4I3776/O  (
    .I(\NlwInverterSignal_MASTER/OE_FRAME/$4I3776/O ),
    .O(\MASTER/OE_FRAME/$4N3742 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$4I3774/I0  (
    .I(OE_AD_T_LT),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$4I3774/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$4I3774/O  (
    .I(\NlwInverterSignal_MASTER/OE_FRAME/$4I3774/O ),
    .O(\MASTER/OE_FRAME/$4N3755 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$4I3772/I0  (
    .I(OE_AD_T_T),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$4I3772/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$4I3772/O  (
    .I(\NlwInverterSignal_MASTER/OE_FRAME/$4I3772/O ),
    .O(\MASTER/OE_FRAME/$4N3754 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$4I3770/I0  (
    .I(\MASTER/OE_FRAME/$4N3742 ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$4I3770/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$4I3770/I1  (
    .I(EOT),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$4I3770/I1 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$4I3770/O  (
    .I(\NlwInverterSignal_MASTER/OE_FRAME/$4I3770/O ),
    .O(\MASTER/OE_FRAME/AD_LB )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$4I3769/I0  (
    .I(\MASTER/OE_FRAME/$4N3755 ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$4I3769/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$4I3769/I1  (
    .I(EOT),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$4I3769/I1 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$4I3769/O  (
    .I(\NlwInverterSignal_MASTER/OE_FRAME/$4I3769/O ),
    .O(\MASTER/OE_FRAME/AD_LT )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$4I3768/I0  (
    .I(\MASTER/OE_FRAME/$4N3754 ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$4I3768/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$4I3768/I1  (
    .I(EOT),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$4I3768/I1 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$4I3768/O  (
    .I(\NlwInverterSignal_MASTER/OE_FRAME/$4I3768/O ),
    .O(\MASTER/OE_FRAME/AD_T )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$3I3105/I0  (
    .I(M_WRDN),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$3I3105/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$3I3105/I1  (
    .I(\MASTER/IIRDY- ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$3I3105/I1 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$3I3105/I2  (
    .I(\TRDY- ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$3I3105/I2 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$3I3105/O  (
    .I(\NlwInverterSignal_MASTER/OE_FRAME/$3I3105/O ),
    .O(\MASTER/OE_FRAME/SET_OE_PERR )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$3I3093/I0  (
    .I(NS_OE_PERR_T),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$3I3093/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$3I3093/I1  (
    .I(\MASTER/OE_FRAME/HOLD_OE_PERR ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$3I3093/I1 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$3I3093/I2  (
    .I(\MASTER/OE_FRAME/SET_OE_PERR ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$3I3093/I2 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$3I3093/O  (
    .I(\NlwInverterSignal_MASTER/OE_FRAME/$3I3093/O ),
    .O(\MASTER/OE_FRAME/NS_OE_PERR )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$2I3723/I0  (
    .I(\GNT- ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$2I3723/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$2I3711/I0  (
    .I(\GNT- ),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$2I3711/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$5I4044/$1I7/I0  (
    .I(SLOT64),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$5I4044/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$5I4044/$1I7/I1  (
    .I(CFG115),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$5I4044/$1I7/I1 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$5I4045/$1I7/I0  (
    .I(SLOT64),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$5I4045/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$5I4045/$1I7/I1  (
    .I(CFG115),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$5I4045/$1I7/I1 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$5I4046/$1I7/I0  (
    .I(SLOT64),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$5I4046/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$5I4046/$1I7/I1  (
    .I(CFG115),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$5I4046/$1I7/I1 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$5I4047/$1I7/I0  (
    .I(SLOT64),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$5I4047/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$5I4047/$1I7/I1  (
    .I(CFG115),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$5I4047/$1I7/I1 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$5I4048/$1I7/I0  (
    .I(SLOT64),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$5I4048/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/OE_FRAME/$5I4048/$1I7/I1  (
    .I(CFG115),
    .O(\NlwInverterSignal_MASTER/OE_FRAME/$5I4048/$1I7/I1 )
  );
  X_INV   \NlwInverterBlock_MASTER/S_TAR/$1I2605/I0  (
    .I(STOP_I),
    .O(\NlwInverterSignal_MASTER/S_TAR/$1I2605/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/DEV_TO/$1I2789/I0  (
    .I(\IFRAME_I- ),
    .O(\NlwInverterSignal_MASTER/DEV_TO/$1I2789/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/DEV_TO/$1I2816/$1I2213/I0  (
    .I(\MASTER/DEV_TO/$1N2820 ),
    .O(\NlwInverterSignal_MASTER/DEV_TO/$1I2816/$1I2213/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/DEV_TO/$1I2838/$1I2213/I0  (
    .I(\MASTER/DEV_TO/$1N2840 ),
    .O(\NlwInverterSignal_MASTER/DEV_TO/$1I2838/$1I2213/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/LAT_TIMR/$2I56/I0  (
    .I(\MASTER/CNT_VAL3 ),
    .O(\NlwInverterSignal_MASTER/LAT_TIMR/$2I56/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/LAT_TIMR/$2I56/I1  (
    .I(\MASTER/CNT_VAL2 ),
    .O(\NlwInverterSignal_MASTER/LAT_TIMR/$2I56/I1 )
  );
  X_INV   \NlwInverterBlock_MASTER/LAT_TIMR/$2I56/I2  (
    .I(\MASTER/CNT_VAL1 ),
    .O(\NlwInverterSignal_MASTER/LAT_TIMR/$2I56/I2 )
  );
  X_INV   \NlwInverterBlock_MASTER/LAT_TIMR/$2I23/I0  (
    .I(\MASTER/CNT_VAL3 ),
    .O(\NlwInverterSignal_MASTER/LAT_TIMR/$2I23/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/LAT_TIMR/$2I23/I1  (
    .I(\MASTER/CNT_VAL2 ),
    .O(\NlwInverterSignal_MASTER/LAT_TIMR/$2I23/I1 )
  );
  X_INV   \NlwInverterBlock_MASTER/LAT_TIMR/$2I23/I2  (
    .I(\MASTER/CNT_VAL1 ),
    .O(\NlwInverterSignal_MASTER/LAT_TIMR/$2I23/I2 )
  );
  X_INV   \NlwInverterBlock_MASTER/LAT_TIMR/$2I23/I3  (
    .I(\MASTER/CNT_VAL0 ),
    .O(\NlwInverterSignal_MASTER/LAT_TIMR/$2I23/I3 )
  );
  X_INV   \NlwInverterBlock_MASTER/LAT_TIMR/$2I21/I0  (
    .I(\MASTER/CNT_VAL2 ),
    .O(\NlwInverterSignal_MASTER/LAT_TIMR/$2I21/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/LAT_TIMR/$2I21/I1  (
    .I(\MASTER/CNT_VAL1 ),
    .O(\NlwInverterSignal_MASTER/LAT_TIMR/$2I21/I1 )
  );
  X_INV   \NlwInverterBlock_MASTER/LAT_TIMR/$2I21/I2  (
    .I(\MASTER/CNT_VAL0 ),
    .O(\NlwInverterSignal_MASTER/LAT_TIMR/$2I21/I2 )
  );
  X_INV   \NlwInverterBlock_MASTER/LAT_TIMR/$2I19/I0  (
    .I(\MASTER/CNT_VAL1 ),
    .O(\NlwInverterSignal_MASTER/LAT_TIMR/$2I19/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/LAT_TIMR/$2I19/I1  (
    .I(\MASTER/CNT_VAL0 ),
    .O(\NlwInverterSignal_MASTER/LAT_TIMR/$2I19/I1 )
  );
  X_INV   \NlwInverterBlock_MASTER/LAT_TIMR/$1I8/I0  (
    .I(\MASTER/CNT_VAL5 ),
    .O(\NlwInverterSignal_MASTER/LAT_TIMR/$1I8/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/LAT_TIMR/$1I8/I1  (
    .I(\MASTER/CNT_VAL4 ),
    .O(\NlwInverterSignal_MASTER/LAT_TIMR/$1I8/I1 )
  );
  X_INV   \NlwInverterBlock_MASTER/LAT_TIMR/$1I29/I0  (
    .I(\MASTER/CNT_VAL7 ),
    .O(\NlwInverterSignal_MASTER/LAT_TIMR/$1I29/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/LAT_TIMR/$1I29/I1  (
    .I(\MASTER/CNT_VAL6 ),
    .O(\NlwInverterSignal_MASTER/LAT_TIMR/$1I29/I1 )
  );
  X_INV   \NlwInverterBlock_MASTER/LAT_TIMR/$1I29/I2  (
    .I(\MASTER/CNT_VAL5 ),
    .O(\NlwInverterSignal_MASTER/LAT_TIMR/$1I29/I2 )
  );
  X_INV   \NlwInverterBlock_MASTER/LAT_TIMR/$1I29/I3  (
    .I(\MASTER/CNT_VAL4 ),
    .O(\NlwInverterSignal_MASTER/LAT_TIMR/$1I29/I3 )
  );
  X_INV   \NlwInverterBlock_MASTER/LAT_TIMR/$1I25/I0  (
    .I(\MASTER/CNT_VAL6 ),
    .O(\NlwInverterSignal_MASTER/LAT_TIMR/$1I25/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/LAT_TIMR/$1I25/I1  (
    .I(\MASTER/CNT_VAL5 ),
    .O(\NlwInverterSignal_MASTER/LAT_TIMR/$1I25/I1 )
  );
  X_INV   \NlwInverterBlock_MASTER/LAT_TIMR/$1I25/I2  (
    .I(\MASTER/CNT_VAL4 ),
    .O(\NlwInverterSignal_MASTER/LAT_TIMR/$1I25/I2 )
  );
  X_INV   \NlwInverterBlock_MASTER/LAT_TIMR/$1I11/I0  (
    .I(\MASTER/CNT_VAL4 ),
    .O(\NlwInverterSignal_MASTER/LAT_TIMR/$1I11/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/LAT_TIMR/Q4/$1I30/$1I7/I0  (
    .I(\IFRAME_I- ),
    .O(\NlwInverterSignal_MASTER/LAT_TIMR/Q4/$1I30/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/LAT_TIMR/Q6/$1I30/$1I7/I0  (
    .I(\IFRAME_I- ),
    .O(\NlwInverterSignal_MASTER/LAT_TIMR/Q6/$1I30/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/LAT_TIMR/Q7/$1I30/$1I7/I0  (
    .I(\IFRAME_I- ),
    .O(\NlwInverterSignal_MASTER/LAT_TIMR/Q7/$1I30/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/LAT_TIMR/TIME_OUT/$1I2214/I0  (
    .I(\MASTER/LAT_TIMR/$1N76 ),
    .O(\NlwInverterSignal_MASTER/LAT_TIMR/TIME_OUT/$1I2214/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/LAT_TIMR/Q5/$1I30/$1I7/I0  (
    .I(\IFRAME_I- ),
    .O(\NlwInverterSignal_MASTER/LAT_TIMR/Q5/$1I30/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/LAT_TIMR/Q1/$1I30/$1I7/I0  (
    .I(\IFRAME_I- ),
    .O(\NlwInverterSignal_MASTER/LAT_TIMR/Q1/$1I30/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/LAT_TIMR/Q0/$1I30/$1I7/I0  (
    .I(\IFRAME_I- ),
    .O(\NlwInverterSignal_MASTER/LAT_TIMR/Q0/$1I30/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/LAT_TIMR/Q2/$1I30/$1I7/I0  (
    .I(\IFRAME_I- ),
    .O(\NlwInverterSignal_MASTER/LAT_TIMR/Q2/$1I30/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/LAT_TIMR/Q3/$1I30/$1I7/I0  (
    .I(\IFRAME_I- ),
    .O(\NlwInverterSignal_MASTER/LAT_TIMR/Q3/$1I30/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_MASTER/3/UPPER/T0/T  (
    .I(OE3),
    .O(\NlwInverterSignal_MASTER/3/UPPER/T0/T )
  );
  X_INV   \NlwInverterBlock_MASTER/3/UPPER/T1/T  (
    .I(OE3),
    .O(\NlwInverterSignal_MASTER/3/UPPER/T1/T )
  );
  X_INV   \NlwInverterBlock_MASTER/3/UPPER/T2/T  (
    .I(OE3),
    .O(\NlwInverterSignal_MASTER/3/UPPER/T2/T )
  );
  X_INV   \NlwInverterBlock_MASTER/3/UPPER/T3/T  (
    .I(OE3),
    .O(\NlwInverterSignal_MASTER/3/UPPER/T3/T )
  );
  X_INV   \NlwInverterBlock_MASTER/3/UPPER/T4/T  (
    .I(OE3),
    .O(\NlwInverterSignal_MASTER/3/UPPER/T4/T )
  );
  X_INV   \NlwInverterBlock_MASTER/3/UPPER/T5/T  (
    .I(OE3),
    .O(\NlwInverterSignal_MASTER/3/UPPER/T5/T )
  );
  X_INV   \NlwInverterBlock_MASTER/3/UPPER/T6/T  (
    .I(OE3),
    .O(\NlwInverterSignal_MASTER/3/UPPER/T6/T )
  );
  X_INV   \NlwInverterBlock_MASTER/3/UPPER/T7/T  (
    .I(OE3),
    .O(\NlwInverterSignal_MASTER/3/UPPER/T7/T )
  );
  X_INV   \NlwInverterBlock_MASTER/3/UPPER/T8/T  (
    .I(OE3),
    .O(\NlwInverterSignal_MASTER/3/UPPER/T8/T )
  );
  X_INV   \NlwInverterBlock_MASTER/3/UPPER/T9/T  (
    .I(OE3),
    .O(\NlwInverterSignal_MASTER/3/UPPER/T9/T )
  );
  X_INV   \NlwInverterBlock_MASTER/3/UPPER/T10/T  (
    .I(OE3),
    .O(\NlwInverterSignal_MASTER/3/UPPER/T10/T )
  );
  X_INV   \NlwInverterBlock_MASTER/3/UPPER/T11/T  (
    .I(OE3),
    .O(\NlwInverterSignal_MASTER/3/UPPER/T11/T )
  );
  X_INV   \NlwInverterBlock_MASTER/3/UPPER/T12/T  (
    .I(OE3),
    .O(\NlwInverterSignal_MASTER/3/UPPER/T12/T )
  );
  X_INV   \NlwInverterBlock_MASTER/3/UPPER/T13/T  (
    .I(OE3),
    .O(\NlwInverterSignal_MASTER/3/UPPER/T13/T )
  );
  X_INV   \NlwInverterBlock_MASTER/3/UPPER/T14/T  (
    .I(OE3),
    .O(\NlwInverterSignal_MASTER/3/UPPER/T14/T )
  );
  X_INV   \NlwInverterBlock_MASTER/3/UPPER/T15/T  (
    .I(OE3),
    .O(\NlwInverterSignal_MASTER/3/UPPER/T15/T )
  );
  X_INV   \NlwInverterBlock_MASTER/3/LOWER/T0/T  (
    .I(OE3),
    .O(\NlwInverterSignal_MASTER/3/LOWER/T0/T )
  );
  X_INV   \NlwInverterBlock_MASTER/3/LOWER/T1/T  (
    .I(OE3),
    .O(\NlwInverterSignal_MASTER/3/LOWER/T1/T )
  );
  X_INV   \NlwInverterBlock_MASTER/3/LOWER/T2/T  (
    .I(OE3),
    .O(\NlwInverterSignal_MASTER/3/LOWER/T2/T )
  );
  X_INV   \NlwInverterBlock_MASTER/3/LOWER/T3/T  (
    .I(OE3),
    .O(\NlwInverterSignal_MASTER/3/LOWER/T3/T )
  );
  X_INV   \NlwInverterBlock_MASTER/3/LOWER/T4/T  (
    .I(OE3),
    .O(\NlwInverterSignal_MASTER/3/LOWER/T4/T )
  );
  X_INV   \NlwInverterBlock_MASTER/3/LOWER/T5/T  (
    .I(OE3),
    .O(\NlwInverterSignal_MASTER/3/LOWER/T5/T )
  );
  X_INV   \NlwInverterBlock_MASTER/3/LOWER/T6/T  (
    .I(OE3),
    .O(\NlwInverterSignal_MASTER/3/LOWER/T6/T )
  );
  X_INV   \NlwInverterBlock_MASTER/3/LOWER/T7/T  (
    .I(OE3),
    .O(\NlwInverterSignal_MASTER/3/LOWER/T7/T )
  );
  X_INV   \NlwInverterBlock_MASTER/3/LOWER/T8/T  (
    .I(OE3),
    .O(\NlwInverterSignal_MASTER/3/LOWER/T8/T )
  );
  X_INV   \NlwInverterBlock_MASTER/3/LOWER/T9/T  (
    .I(OE3),
    .O(\NlwInverterSignal_MASTER/3/LOWER/T9/T )
  );
  X_INV   \NlwInverterBlock_MASTER/3/LOWER/T10/T  (
    .I(OE3),
    .O(\NlwInverterSignal_MASTER/3/LOWER/T10/T )
  );
  X_INV   \NlwInverterBlock_MASTER/3/LOWER/T11/T  (
    .I(OE3),
    .O(\NlwInverterSignal_MASTER/3/LOWER/T11/T )
  );
  X_INV   \NlwInverterBlock_MASTER/3/LOWER/T12/T  (
    .I(OE3),
    .O(\NlwInverterSignal_MASTER/3/LOWER/T12/T )
  );
  X_INV   \NlwInverterBlock_MASTER/3/LOWER/T13/T  (
    .I(OE3),
    .O(\NlwInverterSignal_MASTER/3/LOWER/T13/T )
  );
  X_INV   \NlwInverterBlock_MASTER/3/LOWER/T14/T  (
    .I(OE3),
    .O(\NlwInverterSignal_MASTER/3/LOWER/T14/T )
  );
  X_INV   \NlwInverterBlock_MASTER/3/LOWER/T15/T  (
    .I(OE3),
    .O(\NlwInverterSignal_MASTER/3/LOWER/T15/T )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/$4I788/I0  (
    .I(\TTRDY_I- ),
    .O(\NlwInverterSignal_PCI-CNTL/$4I788/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/$4I719/I0  (
    .I(IRDY_M),
    .O(\NlwInverterSignal_PCI-CNTL/$4I719/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/$4I446/I0  (
    .I(IRDY_M),
    .O(\NlwInverterSignal_PCI-CNTL/$4I446/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/$1I840/I0  (
    .I(\IRDY- ),
    .O(\NlwInverterSignal_PCI-CNTL/$1I840/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/$1I840/I1  (
    .I(\PCI-CNTL/TTRDY- ),
    .O(\NlwInverterSignal_PCI-CNTL/$1I840/I1 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/$1I823/I0  (
    .I(\PCI-CNTL/TDEVSEL- ),
    .O(\NlwInverterSignal_PCI-CNTL/$1I823/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/$1I1005/I0  (
    .I(APERR_N),
    .O(\NlwInverterSignal_PCI-CNTL/$1I1005/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-LC/$2I3201/I0  (
    .I(AD0),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-LC/$2I3201/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-LC/$2I3201/I1  (
    .I(AD1),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-LC/$2I3201/I1 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-LC/$2I3192/I0  (
    .I(CBE_IN2),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-LC/$2I3192/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-LC/$2I3076/I0  (
    .I(IDLE_INT),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-LC/$2I3076/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OE/$2I940/I0  (
    .I(CFG118),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OE/$2I940/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OE/$2I934/I0  (
    .I(CFG0),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OE/$2I934/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OE/$2I933/I0  (
    .I(CFG37),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OE/$2I933/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OE/$2I932/I0  (
    .I(CFG74),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OE/$2I932/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OE/$2I777/I0  (
    .I(NlwRenamedSig_OI_ADDR6),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OE/$2I777/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OE/$2I777/I1  (
    .I(NlwRenamedSig_OI_ADDR7),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OE/$2I777/I1 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OE/$2I592/I0  (
    .I(OLDKEEPOUT),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OE/$2I592/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OE/OE15/$1I307/I0  (
    .I(\PCI-CNTL/PCI-OE/OE15/R ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OE/OE15/$1I307/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OE/OE15/$1I296/I0  (
    .I(OLDKEEPOUT),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OE/OE15/$1I296/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OE/OE7/$1I307/I0  (
    .I(\PCI-CNTL/PCI-OE/OE7/R ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OE/OE7/$1I307/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OE/OE7/$1I296/I0  (
    .I(OLDKEEPOUT),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OE/OE7/$1I296/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OE/OE6/$1I307/I0  (
    .I(\PCI-CNTL/PCI-OE/OE6/R ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OE/OE6/$1I307/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OE/OE6/$1I296/I0  (
    .I(OLDKEEPOUT),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OE/OE6/$1I296/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OE/OE5/$1I307/I0  (
    .I(\PCI-CNTL/PCI-OE/OE5/R ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OE/OE5/$1I307/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OE/OE5/$1I296/I0  (
    .I(OLDKEEPOUT),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OE/OE5/$1I296/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OE/OE4/$1I307/I0  (
    .I(\PCI-CNTL/PCI-OE/OE4/R ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OE/OE4/$1I307/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OE/OE4/$1I296/I0  (
    .I(OLDKEEPOUT),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OE/OE4/$1I296/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OE/OE3/$1I307/I0  (
    .I(\PCI-CNTL/PCI-OE/OE3/R ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OE/OE3/$1I307/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OE/OE3/$1I296/I0  (
    .I(OLDKEEPOUT),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OE/OE3/$1I296/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OE/OE8/$1I307/I0  (
    .I(\PCI-CNTL/PCI-OE/OE8/R ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OE/OE8/$1I307/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OE/OE8/$1I296/I0  (
    .I(OLDKEEPOUT),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OE/OE8/$1I296/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OE/OE9/$1I307/I0  (
    .I(\PCI-CNTL/PCI-OE/OE9/R ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OE/OE9/$1I307/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OE/OE9/$1I296/I0  (
    .I(OLDKEEPOUT),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OE/OE9/$1I296/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OE/OE12/$1I307/I0  (
    .I(\PCI-CNTL/PCI-OE/OE12/R ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OE/OE12/$1I307/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OE/OE12/$1I296/I0  (
    .I(OLDKEEPOUT),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OE/OE12/$1I296/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OE/OE1/$1I307/I0  (
    .I(\PCI-CNTL/PCI-OE/OE1/R ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OE/OE1/$1I307/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OE/OE1/$1I296/I0  (
    .I(OLDKEEPOUT),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OE/OE1/$1I296/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OE/$2I617/$1I11/I0  (
    .I(\PCI-CNTL/PCI-OE/NS_OE_ROM ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OE/$2I617/$1I11/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/$1I995/$1I2213/I0  (
    .I(IDLE_INT),
    .O(\NlwInverterSignal_PCI-CNTL/$1I995/$1I2213/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-TSM/PCI-IDLE/$1I494/I0  (
    .I(\PCI-CNTL/TSTOP- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-IDLE/$1I494/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-TSM/PCI-IDLE/$1I494/I1  (
    .I(\PCI-CNTL/TTRDY- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-IDLE/$1I494/I1 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-TSM/PCI-BUSY/$1I542/I0  (
    .I(\PCI-CNTL/PCI-TSM/PCI-BUSY/HITIDLEORBUSY ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-BUSY/$1I542/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-TSM/PCI-BUSY/$1I521/I0  (
    .I(\PCI-CNTL/PCI-TSM/PCI-BUSY/HITIDLEORBUSY ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-BUSY/$1I521/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-TSM/PCI-BUSY/$1I471/I0  (
    .I(\IRDY- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-BUSY/$1I471/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-TSM/PCI-BUSY/$1I471/I1  (
    .I(\FRAME- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-BUSY/$1I471/I1 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-TSM/PCI-BUSY/$1I469/I0  (
    .I(\FRAME- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-BUSY/$1I469/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-TSM/PCI-DATA/$1I670/I0  (
    .I(\IRDY- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-DATA/$1I670/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-TSM/PCI-DATA/$1I670/I1  (
    .I(\FRAME- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-DATA/$1I670/I1 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-TSM/PCI-DATA/$1I627/I0  (
    .I(C_TERM),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-DATA/$1I627/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-TSM/PCI-DATA/$1I481/I0  (
    .I(\FRAME- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-DATA/$1I481/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-TSM/PCI-DATA/$1I480/I0  (
    .I(\FRAME- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-DATA/$1I480/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-TSM/PCI-DATA/$1I480/I1  (
    .I(\PCI-CNTL/TSTOP- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-DATA/$1I480/I1 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-TSM/PCI-DATA/$1I480/I2  (
    .I(\PCI-CNTL/TTRDY- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-DATA/$1I480/I2 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-TSM/PCI-DATA/$1I453/I0  (
    .I(S_TERM),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-DATA/$1I453/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-TSM/PCI-BKOF/$1I579/I0  (
    .I(S_READY),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-BKOF/$1I579/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-TSM/PCI-BKOF/$1I575/I0  (
    .I(C_READY),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-BKOF/$1I575/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-TSM/PCI-BKOF/$1I526/I0  (
    .I(\IRDY- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-BKOF/$1I526/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-TSM/PCI-BKOF/$1I526/I1  (
    .I(\FRAME- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-BKOF/$1I526/I1 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-TSM/PCI-BKOF/$1I486/I0  (
    .I(\FRAME- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-BKOF/$1I486/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-TSM/PCI-BKOF/$1I475/I0  (
    .I(\IRDY- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-BKOF/$1I475/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-TSM/PCI-BKOF/$1I474/I0  (
    .I(\PCI-CNTL/TSTOP- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-BKOF/$1I474/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-TSM/PCI-BKOF/$1I474/I1  (
    .I(\FRAME- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-BKOF/$1I474/I1 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-TSM/PCI-BKOF/$1I458/I0  (
    .I(\FRAME- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-TSM/PCI-BKOF/$1I458/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-AK64/$3I855/O  (
    .I(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-AK64/$3I855/O ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-AK64/NS_F0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-AK64/$2I971/I0  (
    .I(\PCI-CNTL/S_ABORT ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-AK64/$2I971/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-AK64/$2I965/I0  (
    .I(\PCI-CNTL/PCI-OFCN/PCI-AK64/DUCKLING ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-AK64/$2I965/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-AK64/$2I958/I0  (
    .I(\REQ64- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-AK64/$2I958/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-AK64/$2I951/I0  (
    .I(\REQ64- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-AK64/$2I951/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-AK64/$2I941/I0  (
    .I(\REQ64- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-AK64/$2I941/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-AK64/$1I837/I0  (
    .I(\PCI-CNTL/S_ABORT ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-AK64/$1I837/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-AK64/$1I797/I0  (
    .I(\REQ64- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-AK64/$1I797/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-AK64/$1I796/I0  (
    .I(\REQ64- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-AK64/$1I796/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-AK64/$1I787/O  (
    .I(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-AK64/$1I787/O ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-AK64/NS_F1 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-AK64/$1I781/I0  (
    .I(\IRDY- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-AK64/$1I781/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-AK64/$1I781/I1  (
    .I(\REQ64- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-AK64/$1I781/I1 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-AK64/$3I854/$1I7/I0  (
    .I(IRDY_M),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-AK64/$3I854/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-DSEL/$3I795/O  (
    .I(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-DSEL/$3I795/O ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-DSEL/NS_F0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-DSEL/$2I983/I0  (
    .I(\FRAME- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-DSEL/$2I983/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-DSEL/$2I951/I0  (
    .I(\FRAME- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-DSEL/$2I951/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-DSEL/$2I931/I0  (
    .I(\FRAME- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-DSEL/$2I931/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-DSEL/$2I914/I0  (
    .I(\PCI-CNTL/S_ABORT ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-DSEL/$2I914/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-DSEL/$2I878/I0  (
    .I(\PCI-CNTL/PCI-OFCN/PCI-DSEL/DUCKLING ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-DSEL/$2I878/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-DSEL/$1I801/O  (
    .I(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-DSEL/$1I801/O ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-DSEL/NS_F1 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-DSEL/$1I768/I0  (
    .I(\FRAME- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-DSEL/$1I768/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-DSEL/$1I760/I0  (
    .I(\FRAME- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-DSEL/$1I760/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-DSEL/$1I758/I0  (
    .I(\PCI-CNTL/S_ABORT ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-DSEL/$1I758/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-DSEL/$1I1028/I0  (
    .I(\IRDY- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-DSEL/$1I1028/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-DSEL/$1I1028/I1  (
    .I(\FRAME- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-DSEL/$1I1028/I1 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-DSEL/$3I798/$1I7/I0  (
    .I(IRDY_M),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-DSEL/$3I798/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-TRDY/$4I977/I0  (
    .I(\TSTOP_I- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$4I977/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-TRDY/$4I1044/I0  (
    .I(\TTRDY_I- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$4I1044/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-TRDY/$4I1044/I1  (
    .I(\TSTOP_I- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$4I1044/I1 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-TRDY/$4I1010/I0  (
    .I(\PCI-CNTL/PCI-OFCN/PCI-TRDY/SWAN0 ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$4I1010/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-TRDY/$4I1010/O  (
    .I(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$4I1010/O ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-TRDY/$4N1002 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-TRDY/$3I856/I0  (
    .I(\TTRDY_I- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$3I856/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-TRDY/$3I856/I1  (
    .I(\TSTOP_I- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$3I856/I1 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-TRDY/$3I825/I0  (
    .I(IRDY_M),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$3I825/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-TRDY/$3I823/I0  (
    .I(IRDY_M),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$3I823/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-TRDY/$3I822/I0  (
    .I(\TSTOP_I- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$3I822/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-TRDY/$3I616/I0  (
    .I(\PCI-CNTL/PCI-OFCN/PCI-TRDY/SWAN0 ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$3I616/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-TRDY/$3I616/O  (
    .I(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$3I616/O ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-TRDY/SWAN2 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I785/I0  (
    .I(\PCI-CNTL/S_ABORT ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I785/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I768/I0  (
    .I(\TSTOP_I- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I768/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I746/O  (
    .I(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I746/O ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-TRDY/NS_TRDY- )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I731/I0  (
    .I(C_TERM),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I731/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I481/I0  (
    .I(\FRAME- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I481/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I480/I0  (
    .I(\FRAME- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I480/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I480/I1  (
    .I(\PCI-CNTL/TSTOP- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I480/I1 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I480/I2  (
    .I(\PCI-CNTL/TTRDY- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I480/I2 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I459/I0  (
    .I(\IRDY- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I459/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I459/I1  (
    .I(\FRAME- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I459/I1 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I453/I0  (
    .I(S_TERM),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I453/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I782/$1I7/I0  (
    .I(\PCI-CNTL/CFG_CYC ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$1I782/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-TRDY/$4I1028/$1I7/I0  (
    .I(IRDY_M),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-TRDY/$4I1028/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-STOP/$3I1287/I0  (
    .I(\PCI-CNTL/PCI-OFCN/PCI-STOP/$3N1280 ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$3I1287/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-STOP/$3I1287/O  (
    .I(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$3I1287/O ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-STOP/NS_1 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-STOP/$3I1286/I0  (
    .I(\TSTOP_I- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$3I1286/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-STOP/$3I1284/I0  (
    .I(\TSTOP_I- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$3I1284/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-STOP/$3I1263/I0  (
    .I(\PCI-CNTL/PCI-OFCN/PCI-STOP/$3N1256 ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$3I1263/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-STOP/$3I1263/O  (
    .I(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$3I1263/O ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-STOP/NS_0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-STOP/$3I1260/I0  (
    .I(\TSTOP_I- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$3I1260/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-STOP/$3I1258/I0  (
    .I(\TTRDY_I- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$3I1258/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1504/I0  (
    .I(\PCI-CNTL/PCI-OFCN/PCI-STOP/$1N1503 ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1504/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1480/I0  (
    .I(\PCI-CNTL/PCI-OFCN/PCI-STOP/I_DATA_FLAG ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1480/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1450/I0  (
    .I(\TSTOP_I- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1450/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1248/I0  (
    .I(\PCI-CNTL/S_ABORT ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1248/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1060/I0  (
    .I(\PCI-CNTL/PCI-OFCN/PCI-STOP/READY ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1060/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1368/$1I7/I0  (
    .I(\PCI-CNTL/CFG_CYC ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1368/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1373/$1I7/I0  (
    .I(\PCI-CNTL/CFG_CYC ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1373/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1437/$1I2213/I0  (
    .I(\PCI-CNTL/PCI-OFCN/PCI-STOP/$1N1438 ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1437/$1I2213/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1499/$1I7/I0  (
    .I(\PCI-CNTL/CFG_CYC ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-STOP/$1I1499/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-XOE/$6I970/I0  (
    .I(OE_AD_T_LB64),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$6I970/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-XOE/$6I970/O  (
    .I(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$6I970/O ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/SET_LB64 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-XOE/$6I969/I0  (
    .I(OE_AD_T_LT64),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$6I969/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-XOE/$6I969/O  (
    .I(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$6I969/O ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/SET_LT64 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-XOE/$6I966/I0  (
    .I(OE_AD_T_T64),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$6I966/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-XOE/$6I966/O  (
    .I(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$6I966/O ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/SET_T64 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-XOE/$6I965/I0  (
    .I(OE_AD_T_B64),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$6I965/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-XOE/$6I965/O  (
    .I(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$6I965/O ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/SET_B64 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-XOE/$5I1041/I0  (
    .I(S_TERM),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$5I1041/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-XOE/$5I1035/I0  (
    .I(\TSTOP_I- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$5I1035/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-XOE/$5I1035/I1  (
    .I(\TTRDY_I- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$5I1035/I1 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-XOE/$5I1034/I0  (
    .I(\IRDY- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$5I1034/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-XOE/$5I1034/I1  (
    .I(\FRAME- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$5I1034/I1 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-XOE/$4I909/I0  (
    .I(OE_AD_T_LB),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$4I909/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-XOE/$4I909/O  (
    .I(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$4I909/O ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/SET_LB )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-XOE/$4I908/I0  (
    .I(OE_AD_T_LT),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$4I908/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-XOE/$4I908/O  (
    .I(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$4I908/O ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/SET_LT )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-XOE/$4I905/I0  (
    .I(OE_AD_T_T),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$4I905/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-XOE/$4I905/O  (
    .I(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$4I905/O ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/SET_T )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-XOE/$4I903/I0  (
    .I(OE_AD_T_B),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$4I903/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-XOE/$4I903/O  (
    .I(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$4I903/O ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/SET_B )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-XOE/$3I899/I0  (
    .I(C_TERM),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$3I899/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-XOE/$3I890/I0  (
    .I(\IRDY- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$3I890/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-XOE/$3I890/I1  (
    .I(\FRAME- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$3I890/I1 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-XOE/$3I801/I0  (
    .I(\TSTOP_I- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$3I801/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-XOE/$3I801/I1  (
    .I(\TTRDY_I- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$3I801/I1 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-XOE/$3I627/I0  (
    .I(S_TERM),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$3I627/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-XOE/$2I822/O  (
    .I(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$2I822/O ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/OE_TRDY_IN )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-XOE/$2I1330/I0  (
    .I(\TACK64_I- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$2I1330/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-XOE/$2I1330/I1  (
    .I(\TTRDY_I- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$2I1330/I1 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-XOE/$2I1330/I2  (
    .I(\TSTOP_I- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$2I1330/I2 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-XOE/$2I1265/O  (
    .I(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$2I1265/O ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/OE_ACK64_IN )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-XOE/$2I1014/I0  (
    .I(\TDEVSEL_I- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$2I1014/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-XOE/$2I1014/I1  (
    .I(\TTRDY_I- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$2I1014/I1 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-XOE/$2I1014/I2  (
    .I(\TSTOP_I- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$2I1014/I2 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-XOE/$1I1251/I0  (
    .I(\PCI-CNTL/PCI-OFCN/PCI-XOE/TRDYDEL ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$1I1251/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-XOE/$1I1251/I1  (
    .I(\IRDY- ),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$1I1251/I1 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-XOE/$1I1251/O  (
    .I(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$1I1251/O ),
    .O(\PCI-CNTL/PCI-OFCN/PCI-XOE/SET_OE_PERR )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/PCI-OFCN/PCI-XOE/$1I1247/I0  (
    .I(NlwRenamedSig_OI_PCI_CMD1),
    .O(\NlwInverterSignal_PCI-CNTL/PCI-OFCN/PCI-XOE/$1I1247/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CNTL/$4I614/$1I7/I0  (
    .I(\PCI-CNTL/HOLDCYC ),
    .O(\NlwInverterSignal_PCI-CNTL/$4I614/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_TDLY/$1I315/M01/$1I31/I0  (
    .I(CFG245),
    .O(\NlwInverterSignal_TDLY/$1I315/M01/$1I31/I0 )
  );
  X_INV   \NlwInverterBlock_TDLY/$1I315/M23/$1I31/I0  (
    .I(CFG245),
    .O(\NlwInverterSignal_TDLY/$1I315/M23/$1I31/I0 )
  );
  X_INV   \NlwInverterBlock_TDLY/$1I328/M01/$1I31/I0  (
    .I(CFG245),
    .O(\NlwInverterSignal_TDLY/$1I328/M01/$1I31/I0 )
  );
  X_INV   \NlwInverterBlock_TDLY/$1I328/M23/$1I31/I0  (
    .I(CFG245),
    .O(\NlwInverterSignal_TDLY/$1I328/M23/$1I31/I0 )
  );
  X_INV   \NlwInverterBlock_IDLY/$1I315/M01/$1I31/I0  (
    .I(CFG245),
    .O(\NlwInverterSignal_IDLY/$1I315/M01/$1I31/I0 )
  );
  X_INV   \NlwInverterBlock_IDLY/$1I315/M23/$1I31/I0  (
    .I(CFG245),
    .O(\NlwInverterSignal_IDLY/$1I315/M23/$1I31/I0 )
  );
  X_INV   \NlwInverterBlock_IDLY/$1I328/M01/$1I31/I0  (
    .I(CFG245),
    .O(\NlwInverterSignal_IDLY/$1I328/M01/$1I31/I0 )
  );
  X_INV   \NlwInverterBlock_IDLY/$1I328/M23/$1I31/I0  (
    .I(CFG245),
    .O(\NlwInverterSignal_IDLY/$1I328/M23/$1I31/I0 )
  );
  X_INV   \NlwInverterBlock_DATA_VLD/$1I426/I0  (
    .I(IRDY_M),
    .O(\NlwInverterSignal_DATA_VLD/$1I426/I0 )
  );
  X_INV   \NlwInverterBlock_DATA_VLD/$1I426/I1  (
    .I(\TTRDY_I- ),
    .O(\NlwInverterSignal_DATA_VLD/$1I426/I1 )
  );
  X_INV   \NlwInverterBlock_DATA_VLD/$1I328/I0  (
    .I(TRDY_M),
    .O(\NlwInverterSignal_DATA_VLD/$1I328/I0 )
  );
  X_INV   \NlwInverterBlock_DATA_VLD/$1I328/I1  (
    .I(\IIRDY_I- ),
    .O(\NlwInverterSignal_DATA_VLD/$1I328/I1 )
  );
  X_INV   \NlwInverterBlock_SRC_EN/$1I742/I0  (
    .I(FAIL64_INT),
    .O(\NlwInverterSignal_SRC_EN/$1I742/I0 )
  );
  X_INV   \NlwInverterBlock_SRC_EN/$1I656/I0  (
    .I(NlwRenamedSig_OI_S_WRDN),
    .O(\NlwInverterSignal_SRC_EN/$1I656/I0 )
  );
  X_INV   \NlwInverterBlock_SRC_EN/$1I615/I0  (
    .I(\IFRAME_I- ),
    .O(\NlwInverterSignal_SRC_EN/$1I615/I0 )
  );
  X_INV   \NlwInverterBlock_SRC_EN/$1I558/I0  (
    .I(\TDEVSEL_I- ),
    .O(\NlwInverterSignal_SRC_EN/$1I558/I0 )
  );
  X_INV   \NlwInverterBlock_OUT_CE/$3I1079/I0  (
    .I(\IIRDY_I- ),
    .O(\NlwInverterSignal_OUT_CE/$3I1079/I0 )
  );
  X_INV   \NlwInverterBlock_OUT_CE/$3I1079/O  (
    .I(\NlwInverterSignal_OUT_CE/$3I1079/O ),
    .O(\OUT_CE/M_OK_N )
  );
  X_INV   \NlwInverterBlock_OUT_CE/$3I1078/I0  (
    .I(\TTRDY_I- ),
    .O(\NlwInverterSignal_OUT_CE/$3I1078/I0 )
  );
  X_INV   \NlwInverterBlock_OUT_CE/$3I1078/O  (
    .I(\NlwInverterSignal_OUT_CE/$3I1078/O ),
    .O(\OUT_CE/S_OK_N )
  );
  X_INV   \NlwInverterBlock_OUT_CE/$3I1062/I0  (
    .I(\IIRDY_I- ),
    .O(\NlwInverterSignal_OUT_CE/$3I1062/I0 )
  );
  X_INV   \NlwInverterBlock_OUT_CE/$3I1062/I1  (
    .I(FAIL64_INT),
    .O(\NlwInverterSignal_OUT_CE/$3I1062/I1 )
  );
  X_INV   \NlwInverterBlock_OUT_CE/$3I1061/I0  (
    .I(\TTRDY_I- ),
    .O(\NlwInverterSignal_OUT_CE/$3I1061/I0 )
  );
  X_INV   \NlwInverterBlock_OUT_CE/$3I1061/I1  (
    .I(FAIL64_INT),
    .O(\NlwInverterSignal_OUT_CE/$3I1061/I1 )
  );
  X_INV   \NlwInverterBlock_OUT_CE/$3I1056/I0  (
    .I(FAIL64_INT),
    .O(\NlwInverterSignal_OUT_CE/$3I1056/I0 )
  );
  X_INV   \NlwInverterBlock_OUT_CE/$2I1086/I0  (
    .I(TRDY_F),
    .O(\NlwInverterSignal_OUT_CE/$2I1086/I0 )
  );
  X_INV   \NlwInverterBlock_OUT_CE/$2I1086/I1  (
    .I(\OUT_CE/M_OK_N ),
    .O(\NlwInverterSignal_OUT_CE/$2I1086/I1 )
  );
  X_INV   \NlwInverterBlock_OUT_CE/$2I1085/I0  (
    .I(TRDY_F),
    .O(\NlwInverterSignal_OUT_CE/$2I1085/I0 )
  );
  X_INV   \NlwInverterBlock_OUT_CE/$2I1085/I1  (
    .I(\OUT_CE/M_OK_N ),
    .O(\NlwInverterSignal_OUT_CE/$2I1085/I1 )
  );
  X_INV   \NlwInverterBlock_OUT_CE/$2I1084/I0  (
    .I(\OUT_CE/$2N1067 ),
    .O(\NlwInverterSignal_OUT_CE/$2I1084/I0 )
  );
  X_INV   \NlwInverterBlock_OUT_CE/$2I1084/I1  (
    .I(\OUT_CE/S_OK_N ),
    .O(\NlwInverterSignal_OUT_CE/$2I1084/I1 )
  );
  X_INV   \NlwInverterBlock_OUT_CE/$2I1083/I0  (
    .I(\OUT_CE/$2N1066 ),
    .O(\NlwInverterSignal_OUT_CE/$2I1083/I0 )
  );
  X_INV   \NlwInverterBlock_OUT_CE/$2I1083/I1  (
    .I(\OUT_CE/S_OK_N ),
    .O(\NlwInverterSignal_OUT_CE/$2I1083/I1 )
  );
  X_INV   \NlwInverterBlock_OUT_CE/$2I1015/I0  (
    .I(TRDY_M),
    .O(\NlwInverterSignal_OUT_CE/$2I1015/I0 )
  );
  X_INV   \NlwInverterBlock_OUT_CE/$2I1015/I1  (
    .I(\OUT_CE/M_OK_N ),
    .O(\NlwInverterSignal_OUT_CE/$2I1015/I1 )
  );
  X_INV   \NlwInverterBlock_OUT_CE/$2I1013/I0  (
    .I(TRDY_M),
    .O(\NlwInverterSignal_OUT_CE/$2I1013/I0 )
  );
  X_INV   \NlwInverterBlock_OUT_CE/$2I1013/I1  (
    .I(\OUT_CE/M_OK_N ),
    .O(\NlwInverterSignal_OUT_CE/$2I1013/I1 )
  );
  X_INV   \NlwInverterBlock_OUT_CE/$2I1012/I0  (
    .I(\OUT_CE/$2N1025 ),
    .O(\NlwInverterSignal_OUT_CE/$2I1012/I0 )
  );
  X_INV   \NlwInverterBlock_OUT_CE/$2I1012/I1  (
    .I(\OUT_CE/S_OK_N ),
    .O(\NlwInverterSignal_OUT_CE/$2I1012/I1 )
  );
  X_INV   \NlwInverterBlock_OUT_CE/$2I1007/I0  (
    .I(\OUT_CE/$2N1024 ),
    .O(\NlwInverterSignal_OUT_CE/$2I1007/I0 )
  );
  X_INV   \NlwInverterBlock_OUT_CE/$2I1007/I1  (
    .I(\OUT_CE/S_OK_N ),
    .O(\NlwInverterSignal_OUT_CE/$2I1007/I1 )
  );
  X_INV   \NlwInverterBlock_OUT_CE/$1I980/I0  (
    .I(IRDY_M),
    .O(\NlwInverterSignal_OUT_CE/$1I980/I0 )
  );
  X_INV   \NlwInverterBlock_OUT_CE/$1I976/I0  (
    .I(IRDY_M),
    .O(\NlwInverterSignal_OUT_CE/$1I976/I0 )
  );
  X_INV   \NlwInverterBlock_OUT_CE/$1I975/I0  (
    .I(\OUT_CE/$1N989 ),
    .O(\NlwInverterSignal_OUT_CE/$1I975/I0 )
  );
  X_INV   \NlwInverterBlock_OUT_CE/$1I972/I0  (
    .I(\OUT_CE/$1N968 ),
    .O(\NlwInverterSignal_OUT_CE/$1I972/I0 )
  );
  X_INV   \NlwInverterBlock_OUT_CE/MAGICBOX/PCI_CE/I0  (
    .I(\OUT_CE/FFA_4285 ),
    .O(\NlwInverterSignal_OUT_CE/MAGICBOX/PCI_CE/I0 )
  );
  X_INV   \NlwInverterBlock_OUT_CE/MAGICBOX/PCI_CE/O  (
    .I(\NlwInverterSignal_OUT_CE/MAGICBOX/PCI_CE/O ),
    .O(\OUT_CE/HARD_CE )
  );
  X_INV   \NlwInverterBlock_OUT_CE/MAGICBOX/I3_NAND_TRDY/I0  (
    .I(\OUT_CE/M_OK_N ),
    .O(\NlwInverterSignal_OUT_CE/MAGICBOX/I3_NAND_TRDY/I0 )
  );
  X_INV   \NlwInverterBlock_OUT_CE/MAGICBOX/I3_NAND_TRDY/I1  (
    .I(TRDY_I),
    .O(\NlwInverterSignal_OUT_CE/MAGICBOX/I3_NAND_TRDY/I1 )
  );
  X_INV   \NlwInverterBlock_OUT_CE/MAGICBOX/I3_NAND_TRDY/O  (
    .I(\NlwInverterSignal_OUT_CE/MAGICBOX/I3_NAND_TRDY/O ),
    .O(\OUT_CE/MAGICBOX/I3_NAND_TRDY_4239 )
  );
  X_INV   \NlwInverterBlock_OUT_CE/MAGICBOX/I1_NAND_IRDY/I0  (
    .I(\OUT_CE/S_OK_N ),
    .O(\NlwInverterSignal_OUT_CE/MAGICBOX/I1_NAND_IRDY/I0 )
  );
  X_INV   \NlwInverterBlock_OUT_CE/MAGICBOX/I1_NAND_IRDY/I1  (
    .I(IRDY_I),
    .O(\NlwInverterSignal_OUT_CE/MAGICBOX/I1_NAND_IRDY/I1 )
  );
  X_INV   \NlwInverterBlock_OUT_CE/MAGICBOX/I1_NAND_IRDY/O  (
    .I(\NlwInverterSignal_OUT_CE/MAGICBOX/I1_NAND_IRDY/O ),
    .O(\OUT_CE/MAGICBOX/I1_NAND_IRDY_4238 )
  );
  X_INV   \NlwInverterBlock_OUT_CE/$4I1005/$1I7/I0  (
    .I(CFG251),
    .O(\NlwInverterSignal_OUT_CE/$4I1005/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_OUT_SEL/$1I916/I0  (
    .I(S_FIRST),
    .O(\NlwInverterSignal_OUT_SEL/$1I916/I0 )
  );
  X_INV   \NlwInverterBlock_OUT_SEL/$1I916/I1  (
    .I(\TDEVSEL_I- ),
    .O(\NlwInverterSignal_OUT_SEL/$1I916/I1 )
  );
  X_INV   \NlwInverterBlock_OUT_SEL/$1I913/I0  (
    .I(ADDR_BE),
    .O(\NlwInverterSignal_OUT_SEL/$1I913/I0 )
  );
  X_INV   \NlwInverterBlock_OUT_SEL/$1I913/I1  (
    .I(M_FIRST),
    .O(\NlwInverterSignal_OUT_SEL/$1I913/I1 )
  );
  X_INV   \NlwInverterBlock_OUT_SEL/$1I913/I2  (
    .I(\IFRAME_I- ),
    .O(\NlwInverterSignal_OUT_SEL/$1I913/I2 )
  );
  X_INV   \NlwInverterBlock_OUT_SEL/$1I897/I0  (
    .I(NlwRenamedSig_OI_S_WRDN),
    .O(\NlwInverterSignal_OUT_SEL/$1I897/I0 )
  );
  X_INV   \NlwInverterBlock_OUT_SEL/$1I853/I0  (
    .I(OUT_SEL64),
    .O(\NlwInverterSignal_OUT_SEL/$1I853/I0 )
  );
  X_INV   \NlwInverterBlock_OUT_SEL/$1I849/I0  (
    .I(OUT_SEL),
    .O(\NlwInverterSignal_OUT_SEL/$1I849/I0 )
  );
  X_INV   \NlwInverterBlock_OUT_SEL/$1I758/I0  (
    .I(NlwRenamedSig_OI_S_WRDN),
    .O(\NlwInverterSignal_OUT_SEL/$1I758/I0 )
  );
  X_INV   \NlwInverterBlock_ADDR_VLD/$1I4008/I0  (
    .I(\REQ64- ),
    .O(\NlwInverterSignal_ADDR_VLD/$1I4008/I0 )
  );
  X_INV   \NlwInverterBlock_ADDR_VLD/$1I4008/I1  (
    .I(\FRAME- ),
    .O(\NlwInverterSignal_ADDR_VLD/$1I4008/I1 )
  );
  X_INV   \NlwInverterBlock_ADDR_VLD/$1I4005/I0  (
    .I(CFG_SELF),
    .O(\NlwInverterSignal_ADDR_VLD/$1I4005/I0 )
  );
  X_INV   \NlwInverterBlock_ADDR_VLD/$1I4005/O  (
    .I(\NlwInverterSignal_ADDR_VLD/$1I4005/O ),
    .O(\ADDR_VLD/TEMP_2 )
  );
  X_INV   \NlwInverterBlock_ADDR_VLD/$1I3989/I0  (
    .I(CFG_SELF),
    .O(\NlwInverterSignal_ADDR_VLD/$1I3989/I0 )
  );
  X_INV   \NlwInverterBlock_ADDR_VLD/$1I3989/O  (
    .I(\NlwInverterSignal_ADDR_VLD/$1I3989/O ),
    .O(\ADDR_VLD/$1N3964 )
  );
  X_INV   \NlwInverterBlock_ADDR_VLD/$1I3986/I0  (
    .I(CFG_SELF),
    .O(\NlwInverterSignal_ADDR_VLD/$1I3986/I0 )
  );
  X_INV   \NlwInverterBlock_ADDR_VLD/$1I3986/O  (
    .I(\NlwInverterSignal_ADDR_VLD/$1I3986/O ),
    .O(\ADDR_VLD/$1N3898 )
  );
  X_INV   \NlwInverterBlock_ADDR_VLD/$1I3983/I0  (
    .I(CFG_SELF),
    .O(\NlwInverterSignal_ADDR_VLD/$1I3983/I0 )
  );
  X_INV   \NlwInverterBlock_ADDR_VLD/$1I3983/O  (
    .I(\NlwInverterSignal_ADDR_VLD/$1I3983/O ),
    .O(\ADDR_VLD/$1N3884 )
  );
  X_INV   \NlwInverterBlock_ADDR_VLD/$1I3980/I0  (
    .I(CFG_SELF),
    .O(\NlwInverterSignal_ADDR_VLD/$1I3980/I0 )
  );
  X_INV   \NlwInverterBlock_ADDR_VLD/$1I3980/O  (
    .I(\NlwInverterSignal_ADDR_VLD/$1I3980/O ),
    .O(\ADDR_VLD/$1N3858 )
  );
  X_INV   \NlwInverterBlock_ADDR_VLD/$1I3963/I0  (
    .I(\FRAME- ),
    .O(\NlwInverterSignal_ADDR_VLD/$1I3963/I0 )
  );
  X_INV   \NlwInverterBlock_ADDR_VLD/$1I3894/I0  (
    .I(\FRAME- ),
    .O(\NlwInverterSignal_ADDR_VLD/$1I3894/I0 )
  );
  X_INV   \NlwInverterBlock_ADDR_VLD/$1I3880/I0  (
    .I(\FRAME- ),
    .O(\NlwInverterSignal_ADDR_VLD/$1I3880/I0 )
  );
  X_INV   \NlwInverterBlock_ADDR_VLD/$1I3867/I0  (
    .I(\FRAME- ),
    .O(\NlwInverterSignal_ADDR_VLD/$1I3867/I0 )
  );
  X_INV   \NlwInverterBlock_EOT/$1I617/I0  (
    .I(STOP_I),
    .O(\NlwInverterSignal_EOT/$1I617/I0 )
  );
  X_INV   \NlwInverterBlock_EOT/$1I617/I1  (
    .I(TRDY_M),
    .O(\NlwInverterSignal_EOT/$1I617/I1 )
  );
  X_INV   \NlwInverterBlock_EOT/$1I616/I0  (
    .I(\EOT/EOT_DL_4369 ),
    .O(\NlwInverterSignal_EOT/$1I616/I0 )
  );
  X_INV   \NlwInverterBlock_EOT/$1I615/I0  (
    .I(\TSTOP_I- ),
    .O(\NlwInverterSignal_EOT/$1I615/I0 )
  );
  X_INV   \NlwInverterBlock_EOT/$1I615/I1  (
    .I(\TTRDY_I- ),
    .O(\NlwInverterSignal_EOT/$1I615/I1 )
  );
  X_INV   \NlwInverterBlock_EOT/$1I589/I0  (
    .I(STOP_I),
    .O(\NlwInverterSignal_EOT/$1I589/I0 )
  );
  X_INV   \NlwInverterBlock_EOT/$1I589/I1  (
    .I(TRDY_M),
    .O(\NlwInverterSignal_EOT/$1I589/I1 )
  );
  X_INV   \NlwInverterBlock_EOT/$1I588/I0  (
    .I(\EOT/EOT_DL_4369 ),
    .O(\NlwInverterSignal_EOT/$1I588/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-PAR/$7I2985/O  (
    .I(\NlwInverterSignal_PCI-PAR/$7I2985/O ),
    .O(\PCI-PAR/PREN )
  );
  X_INV   \NlwInverterBlock_PCI-PAR/$7I2974/O  (
    .I(\NlwInverterSignal_PCI-PAR/$7I2974/O ),
    .O(\PCI-PAR/PRE64N )
  );
  X_INV   \NlwInverterBlock_PCI-PAR/$4I3127/O  (
    .I(\NlwInverterSignal_PCI-PAR/$4I3127/O ),
    .O(\PCI-PAR/PAP_0 )
  );
  X_INV   \NlwInverterBlock_PCI-PAR/$4I3104/O  (
    .I(\NlwInverterSignal_PCI-PAR/$4I3104/O ),
    .O(\PCI-PAR/PAP_1 )
  );
  X_INV   \NlwInverterBlock_PCI-PAR/$3I3057/I0  (
    .I(\PERR- ),
    .O(\NlwInverterSignal_PCI-PAR/$3I3057/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-PAR/$3I3018/O  (
    .I(\NlwInverterSignal_PCI-PAR/$3I3018/O ),
    .O(\PCI-PAR/NS_1 )
  );
  X_INV   \NlwInverterBlock_PCI-PAR/$3I2993/O  (
    .I(\NlwInverterSignal_PCI-PAR/$3I2993/O ),
    .O(\PCI-PAR/NS_0 )
  );
  X_INV   \NlwInverterBlock_PCI-PAR/$3I2940/O  (
    .I(\NlwInverterSignal_PCI-PAR/$3I2940/O ),
    .O(\PCI-PAR/$3N2935 )
  );
  X_INV   \NlwInverterBlock_PCI-PAR/$3I2936/I0  (
    .I(SERR_EN),
    .O(\NlwInverterSignal_PCI-PAR/$3I2936/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-PAR/$3I2931/I0  (
    .I(\PCI-PAR/LC_PERR- ),
    .O(\NlwInverterSignal_PCI-PAR/$3I2931/I0 )
  );
  X_INV   \NlwInverterBlock_4/UPPER/T0/T  (
    .I(BAR0_T),
    .O(\NlwInverterSignal_4/UPPER/T0/T )
  );
  X_INV   \NlwInverterBlock_4/UPPER/T1/T  (
    .I(BAR0_T),
    .O(\NlwInverterSignal_4/UPPER/T1/T )
  );
  X_INV   \NlwInverterBlock_4/UPPER/T2/T  (
    .I(BAR0_T),
    .O(\NlwInverterSignal_4/UPPER/T2/T )
  );
  X_INV   \NlwInverterBlock_4/UPPER/T3/T  (
    .I(BAR0_T),
    .O(\NlwInverterSignal_4/UPPER/T3/T )
  );
  X_INV   \NlwInverterBlock_4/UPPER/T4/T  (
    .I(BAR0_T),
    .O(\NlwInverterSignal_4/UPPER/T4/T )
  );
  X_INV   \NlwInverterBlock_4/UPPER/T5/T  (
    .I(BAR0_T),
    .O(\NlwInverterSignal_4/UPPER/T5/T )
  );
  X_INV   \NlwInverterBlock_4/UPPER/T6/T  (
    .I(BAR0_T),
    .O(\NlwInverterSignal_4/UPPER/T6/T )
  );
  X_INV   \NlwInverterBlock_4/UPPER/T7/T  (
    .I(BAR0_T),
    .O(\NlwInverterSignal_4/UPPER/T7/T )
  );
  X_INV   \NlwInverterBlock_4/UPPER/T8/T  (
    .I(BAR0_T),
    .O(\NlwInverterSignal_4/UPPER/T8/T )
  );
  X_INV   \NlwInverterBlock_4/UPPER/T9/T  (
    .I(BAR0_T),
    .O(\NlwInverterSignal_4/UPPER/T9/T )
  );
  X_INV   \NlwInverterBlock_4/UPPER/T10/T  (
    .I(BAR0_T),
    .O(\NlwInverterSignal_4/UPPER/T10/T )
  );
  X_INV   \NlwInverterBlock_4/UPPER/T11/T  (
    .I(BAR0_T),
    .O(\NlwInverterSignal_4/UPPER/T11/T )
  );
  X_INV   \NlwInverterBlock_4/UPPER/T12/T  (
    .I(BAR0_T),
    .O(\NlwInverterSignal_4/UPPER/T12/T )
  );
  X_INV   \NlwInverterBlock_4/UPPER/T13/T  (
    .I(BAR0_T),
    .O(\NlwInverterSignal_4/UPPER/T13/T )
  );
  X_INV   \NlwInverterBlock_4/UPPER/T14/T  (
    .I(BAR0_T),
    .O(\NlwInverterSignal_4/UPPER/T14/T )
  );
  X_INV   \NlwInverterBlock_4/UPPER/T15/T  (
    .I(BAR0_T),
    .O(\NlwInverterSignal_4/UPPER/T15/T )
  );
  X_INV   \NlwInverterBlock_4/LOWER/T0/T  (
    .I(BAR0_T),
    .O(\NlwInverterSignal_4/LOWER/T0/T )
  );
  X_INV   \NlwInverterBlock_4/LOWER/T1/T  (
    .I(BAR0_T),
    .O(\NlwInverterSignal_4/LOWER/T1/T )
  );
  X_INV   \NlwInverterBlock_4/LOWER/T2/T  (
    .I(BAR0_T),
    .O(\NlwInverterSignal_4/LOWER/T2/T )
  );
  X_INV   \NlwInverterBlock_4/LOWER/T3/T  (
    .I(BAR0_T),
    .O(\NlwInverterSignal_4/LOWER/T3/T )
  );
  X_INV   \NlwInverterBlock_4/LOWER/T4/T  (
    .I(BAR0_T),
    .O(\NlwInverterSignal_4/LOWER/T4/T )
  );
  X_INV   \NlwInverterBlock_4/LOWER/T5/T  (
    .I(BAR0_T),
    .O(\NlwInverterSignal_4/LOWER/T5/T )
  );
  X_INV   \NlwInverterBlock_4/LOWER/T6/T  (
    .I(BAR0_T),
    .O(\NlwInverterSignal_4/LOWER/T6/T )
  );
  X_INV   \NlwInverterBlock_4/LOWER/T7/T  (
    .I(BAR0_T),
    .O(\NlwInverterSignal_4/LOWER/T7/T )
  );
  X_INV   \NlwInverterBlock_4/LOWER/T8/T  (
    .I(BAR0_T),
    .O(\NlwInverterSignal_4/LOWER/T8/T )
  );
  X_INV   \NlwInverterBlock_4/LOWER/T9/T  (
    .I(BAR0_T),
    .O(\NlwInverterSignal_4/LOWER/T9/T )
  );
  X_INV   \NlwInverterBlock_4/LOWER/T10/T  (
    .I(BAR0_T),
    .O(\NlwInverterSignal_4/LOWER/T10/T )
  );
  X_INV   \NlwInverterBlock_4/LOWER/T11/T  (
    .I(BAR0_T),
    .O(\NlwInverterSignal_4/LOWER/T11/T )
  );
  X_INV   \NlwInverterBlock_4/LOWER/T12/T  (
    .I(BAR0_T),
    .O(\NlwInverterSignal_4/LOWER/T12/T )
  );
  X_INV   \NlwInverterBlock_4/LOWER/T13/T  (
    .I(BAR0_T),
    .O(\NlwInverterSignal_4/LOWER/T13/T )
  );
  X_INV   \NlwInverterBlock_4/LOWER/T14/T  (
    .I(BAR0_T),
    .O(\NlwInverterSignal_4/LOWER/T14/T )
  );
  X_INV   \NlwInverterBlock_4/LOWER/T15/T  (
    .I(BAR0_T),
    .O(\NlwInverterSignal_4/LOWER/T15/T )
  );
  X_INV   \NlwInverterBlock_5/UPPER/T0/T  (
    .I(BAR1_T),
    .O(\NlwInverterSignal_5/UPPER/T0/T )
  );
  X_INV   \NlwInverterBlock_5/UPPER/T1/T  (
    .I(BAR1_T),
    .O(\NlwInverterSignal_5/UPPER/T1/T )
  );
  X_INV   \NlwInverterBlock_5/UPPER/T2/T  (
    .I(BAR1_T),
    .O(\NlwInverterSignal_5/UPPER/T2/T )
  );
  X_INV   \NlwInverterBlock_5/UPPER/T3/T  (
    .I(BAR1_T),
    .O(\NlwInverterSignal_5/UPPER/T3/T )
  );
  X_INV   \NlwInverterBlock_5/UPPER/T4/T  (
    .I(BAR1_T),
    .O(\NlwInverterSignal_5/UPPER/T4/T )
  );
  X_INV   \NlwInverterBlock_5/UPPER/T5/T  (
    .I(BAR1_T),
    .O(\NlwInverterSignal_5/UPPER/T5/T )
  );
  X_INV   \NlwInverterBlock_5/UPPER/T6/T  (
    .I(BAR1_T),
    .O(\NlwInverterSignal_5/UPPER/T6/T )
  );
  X_INV   \NlwInverterBlock_5/UPPER/T7/T  (
    .I(BAR1_T),
    .O(\NlwInverterSignal_5/UPPER/T7/T )
  );
  X_INV   \NlwInverterBlock_5/UPPER/T8/T  (
    .I(BAR1_T),
    .O(\NlwInverterSignal_5/UPPER/T8/T )
  );
  X_INV   \NlwInverterBlock_5/UPPER/T9/T  (
    .I(BAR1_T),
    .O(\NlwInverterSignal_5/UPPER/T9/T )
  );
  X_INV   \NlwInverterBlock_5/UPPER/T10/T  (
    .I(BAR1_T),
    .O(\NlwInverterSignal_5/UPPER/T10/T )
  );
  X_INV   \NlwInverterBlock_5/UPPER/T11/T  (
    .I(BAR1_T),
    .O(\NlwInverterSignal_5/UPPER/T11/T )
  );
  X_INV   \NlwInverterBlock_5/UPPER/T12/T  (
    .I(BAR1_T),
    .O(\NlwInverterSignal_5/UPPER/T12/T )
  );
  X_INV   \NlwInverterBlock_5/UPPER/T13/T  (
    .I(BAR1_T),
    .O(\NlwInverterSignal_5/UPPER/T13/T )
  );
  X_INV   \NlwInverterBlock_5/UPPER/T14/T  (
    .I(BAR1_T),
    .O(\NlwInverterSignal_5/UPPER/T14/T )
  );
  X_INV   \NlwInverterBlock_5/UPPER/T15/T  (
    .I(BAR1_T),
    .O(\NlwInverterSignal_5/UPPER/T15/T )
  );
  X_INV   \NlwInverterBlock_5/LOWER/T0/T  (
    .I(BAR1_T),
    .O(\NlwInverterSignal_5/LOWER/T0/T )
  );
  X_INV   \NlwInverterBlock_5/LOWER/T1/T  (
    .I(BAR1_T),
    .O(\NlwInverterSignal_5/LOWER/T1/T )
  );
  X_INV   \NlwInverterBlock_5/LOWER/T2/T  (
    .I(BAR1_T),
    .O(\NlwInverterSignal_5/LOWER/T2/T )
  );
  X_INV   \NlwInverterBlock_5/LOWER/T3/T  (
    .I(BAR1_T),
    .O(\NlwInverterSignal_5/LOWER/T3/T )
  );
  X_INV   \NlwInverterBlock_5/LOWER/T4/T  (
    .I(BAR1_T),
    .O(\NlwInverterSignal_5/LOWER/T4/T )
  );
  X_INV   \NlwInverterBlock_5/LOWER/T5/T  (
    .I(BAR1_T),
    .O(\NlwInverterSignal_5/LOWER/T5/T )
  );
  X_INV   \NlwInverterBlock_5/LOWER/T6/T  (
    .I(BAR1_T),
    .O(\NlwInverterSignal_5/LOWER/T6/T )
  );
  X_INV   \NlwInverterBlock_5/LOWER/T7/T  (
    .I(BAR1_T),
    .O(\NlwInverterSignal_5/LOWER/T7/T )
  );
  X_INV   \NlwInverterBlock_5/LOWER/T8/T  (
    .I(BAR1_T),
    .O(\NlwInverterSignal_5/LOWER/T8/T )
  );
  X_INV   \NlwInverterBlock_5/LOWER/T9/T  (
    .I(BAR1_T),
    .O(\NlwInverterSignal_5/LOWER/T9/T )
  );
  X_INV   \NlwInverterBlock_5/LOWER/T10/T  (
    .I(BAR1_T),
    .O(\NlwInverterSignal_5/LOWER/T10/T )
  );
  X_INV   \NlwInverterBlock_5/LOWER/T11/T  (
    .I(BAR1_T),
    .O(\NlwInverterSignal_5/LOWER/T11/T )
  );
  X_INV   \NlwInverterBlock_5/LOWER/T12/T  (
    .I(BAR1_T),
    .O(\NlwInverterSignal_5/LOWER/T12/T )
  );
  X_INV   \NlwInverterBlock_5/LOWER/T13/T  (
    .I(BAR1_T),
    .O(\NlwInverterSignal_5/LOWER/T13/T )
  );
  X_INV   \NlwInverterBlock_5/LOWER/T14/T  (
    .I(BAR1_T),
    .O(\NlwInverterSignal_5/LOWER/T14/T )
  );
  X_INV   \NlwInverterBlock_5/LOWER/T15/T  (
    .I(BAR1_T),
    .O(\NlwInverterSignal_5/LOWER/T15/T )
  );
  X_INV   \NlwInverterBlock_6/UPPER/T0/T  (
    .I(BAR2_T),
    .O(\NlwInverterSignal_6/UPPER/T0/T )
  );
  X_INV   \NlwInverterBlock_6/UPPER/T1/T  (
    .I(BAR2_T),
    .O(\NlwInverterSignal_6/UPPER/T1/T )
  );
  X_INV   \NlwInverterBlock_6/UPPER/T2/T  (
    .I(BAR2_T),
    .O(\NlwInverterSignal_6/UPPER/T2/T )
  );
  X_INV   \NlwInverterBlock_6/UPPER/T3/T  (
    .I(BAR2_T),
    .O(\NlwInverterSignal_6/UPPER/T3/T )
  );
  X_INV   \NlwInverterBlock_6/UPPER/T4/T  (
    .I(BAR2_T),
    .O(\NlwInverterSignal_6/UPPER/T4/T )
  );
  X_INV   \NlwInverterBlock_6/UPPER/T5/T  (
    .I(BAR2_T),
    .O(\NlwInverterSignal_6/UPPER/T5/T )
  );
  X_INV   \NlwInverterBlock_6/UPPER/T6/T  (
    .I(BAR2_T),
    .O(\NlwInverterSignal_6/UPPER/T6/T )
  );
  X_INV   \NlwInverterBlock_6/UPPER/T7/T  (
    .I(BAR2_T),
    .O(\NlwInverterSignal_6/UPPER/T7/T )
  );
  X_INV   \NlwInverterBlock_6/UPPER/T8/T  (
    .I(BAR2_T),
    .O(\NlwInverterSignal_6/UPPER/T8/T )
  );
  X_INV   \NlwInverterBlock_6/UPPER/T9/T  (
    .I(BAR2_T),
    .O(\NlwInverterSignal_6/UPPER/T9/T )
  );
  X_INV   \NlwInverterBlock_6/UPPER/T10/T  (
    .I(BAR2_T),
    .O(\NlwInverterSignal_6/UPPER/T10/T )
  );
  X_INV   \NlwInverterBlock_6/UPPER/T11/T  (
    .I(BAR2_T),
    .O(\NlwInverterSignal_6/UPPER/T11/T )
  );
  X_INV   \NlwInverterBlock_6/UPPER/T12/T  (
    .I(BAR2_T),
    .O(\NlwInverterSignal_6/UPPER/T12/T )
  );
  X_INV   \NlwInverterBlock_6/UPPER/T13/T  (
    .I(BAR2_T),
    .O(\NlwInverterSignal_6/UPPER/T13/T )
  );
  X_INV   \NlwInverterBlock_6/UPPER/T14/T  (
    .I(BAR2_T),
    .O(\NlwInverterSignal_6/UPPER/T14/T )
  );
  X_INV   \NlwInverterBlock_6/UPPER/T15/T  (
    .I(BAR2_T),
    .O(\NlwInverterSignal_6/UPPER/T15/T )
  );
  X_INV   \NlwInverterBlock_6/LOWER/T0/T  (
    .I(BAR2_T),
    .O(\NlwInverterSignal_6/LOWER/T0/T )
  );
  X_INV   \NlwInverterBlock_6/LOWER/T1/T  (
    .I(BAR2_T),
    .O(\NlwInverterSignal_6/LOWER/T1/T )
  );
  X_INV   \NlwInverterBlock_6/LOWER/T2/T  (
    .I(BAR2_T),
    .O(\NlwInverterSignal_6/LOWER/T2/T )
  );
  X_INV   \NlwInverterBlock_6/LOWER/T3/T  (
    .I(BAR2_T),
    .O(\NlwInverterSignal_6/LOWER/T3/T )
  );
  X_INV   \NlwInverterBlock_6/LOWER/T4/T  (
    .I(BAR2_T),
    .O(\NlwInverterSignal_6/LOWER/T4/T )
  );
  X_INV   \NlwInverterBlock_6/LOWER/T5/T  (
    .I(BAR2_T),
    .O(\NlwInverterSignal_6/LOWER/T5/T )
  );
  X_INV   \NlwInverterBlock_6/LOWER/T6/T  (
    .I(BAR2_T),
    .O(\NlwInverterSignal_6/LOWER/T6/T )
  );
  X_INV   \NlwInverterBlock_6/LOWER/T7/T  (
    .I(BAR2_T),
    .O(\NlwInverterSignal_6/LOWER/T7/T )
  );
  X_INV   \NlwInverterBlock_6/LOWER/T8/T  (
    .I(BAR2_T),
    .O(\NlwInverterSignal_6/LOWER/T8/T )
  );
  X_INV   \NlwInverterBlock_6/LOWER/T9/T  (
    .I(BAR2_T),
    .O(\NlwInverterSignal_6/LOWER/T9/T )
  );
  X_INV   \NlwInverterBlock_6/LOWER/T10/T  (
    .I(BAR2_T),
    .O(\NlwInverterSignal_6/LOWER/T10/T )
  );
  X_INV   \NlwInverterBlock_6/LOWER/T11/T  (
    .I(BAR2_T),
    .O(\NlwInverterSignal_6/LOWER/T11/T )
  );
  X_INV   \NlwInverterBlock_6/LOWER/T12/T  (
    .I(BAR2_T),
    .O(\NlwInverterSignal_6/LOWER/T12/T )
  );
  X_INV   \NlwInverterBlock_6/LOWER/T13/T  (
    .I(BAR2_T),
    .O(\NlwInverterSignal_6/LOWER/T13/T )
  );
  X_INV   \NlwInverterBlock_6/LOWER/T14/T  (
    .I(BAR2_T),
    .O(\NlwInverterSignal_6/LOWER/T14/T )
  );
  X_INV   \NlwInverterBlock_6/LOWER/T15/T  (
    .I(BAR2_T),
    .O(\NlwInverterSignal_6/LOWER/T15/T )
  );
  X_INV   \NlwInverterBlock_BAR0/BR-31-24/X1/O  (
    .I(\NlwInverterSignal_BAR0/BR-31-24/X1/O ),
    .O(\BAR0/BR-31-24/EQ1 )
  );
  X_INV   \NlwInverterBlock_BAR0/BR-31-24/X3/O  (
    .I(\NlwInverterSignal_BAR0/BR-31-24/X3/O ),
    .O(\BAR0/BR-31-24/EQ3 )
  );
  X_INV   \NlwInverterBlock_BAR0/BR-31-24/X2/O  (
    .I(\NlwInverterSignal_BAR0/BR-31-24/X2/O ),
    .O(\BAR0/BR-31-24/EQ2 )
  );
  X_INV   \NlwInverterBlock_BAR0/BR-31-24/X0/O  (
    .I(\NlwInverterSignal_BAR0/BR-31-24/X0/O ),
    .O(\BAR0/BR-31-24/EQ0 )
  );
  X_INV   \NlwInverterBlock_BAR0/BR-31-24/X4/O  (
    .I(\NlwInverterSignal_BAR0/BR-31-24/X4/O ),
    .O(\BAR0/BR-31-24/EQ4 )
  );
  X_INV   \NlwInverterBlock_BAR0/BR-31-24/X6/O  (
    .I(\NlwInverterSignal_BAR0/BR-31-24/X6/O ),
    .O(\BAR0/BR-31-24/EQ6 )
  );
  X_INV   \NlwInverterBlock_BAR0/BR-31-24/X7/O  (
    .I(\NlwInverterSignal_BAR0/BR-31-24/X7/O ),
    .O(\BAR0/BR-31-24/EQ7 )
  );
  X_INV   \NlwInverterBlock_BAR0/BR-31-24/X5/O  (
    .I(\NlwInverterSignal_BAR0/BR-31-24/X5/O ),
    .O(\BAR0/BR-31-24/EQ5 )
  );
  X_INV   \NlwInverterBlock_BAR0/BR-23-16/X1/O  (
    .I(\NlwInverterSignal_BAR0/BR-23-16/X1/O ),
    .O(\BAR0/BR-23-16/EQ1 )
  );
  X_INV   \NlwInverterBlock_BAR0/BR-23-16/X3/O  (
    .I(\NlwInverterSignal_BAR0/BR-23-16/X3/O ),
    .O(\BAR0/BR-23-16/EQ3 )
  );
  X_INV   \NlwInverterBlock_BAR0/BR-23-16/X2/O  (
    .I(\NlwInverterSignal_BAR0/BR-23-16/X2/O ),
    .O(\BAR0/BR-23-16/EQ2 )
  );
  X_INV   \NlwInverterBlock_BAR0/BR-23-16/X0/O  (
    .I(\NlwInverterSignal_BAR0/BR-23-16/X0/O ),
    .O(\BAR0/BR-23-16/EQ0 )
  );
  X_INV   \NlwInverterBlock_BAR0/BR-23-16/X4/O  (
    .I(\NlwInverterSignal_BAR0/BR-23-16/X4/O ),
    .O(\BAR0/BR-23-16/EQ4 )
  );
  X_INV   \NlwInverterBlock_BAR0/BR-23-16/X6/O  (
    .I(\NlwInverterSignal_BAR0/BR-23-16/X6/O ),
    .O(\BAR0/BR-23-16/EQ6 )
  );
  X_INV   \NlwInverterBlock_BAR0/BR-23-16/X7/O  (
    .I(\NlwInverterSignal_BAR0/BR-23-16/X7/O ),
    .O(\BAR0/BR-23-16/EQ7 )
  );
  X_INV   \NlwInverterBlock_BAR0/BR-23-16/X5/O  (
    .I(\NlwInverterSignal_BAR0/BR-23-16/X5/O ),
    .O(\BAR0/BR-23-16/EQ5 )
  );
  X_INV   \NlwInverterBlock_BAR0/BR-15-8/X1/O  (
    .I(\NlwInverterSignal_BAR0/BR-15-8/X1/O ),
    .O(\BAR0/BR-15-8/EQ1 )
  );
  X_INV   \NlwInverterBlock_BAR0/BR-15-8/X3/O  (
    .I(\NlwInverterSignal_BAR0/BR-15-8/X3/O ),
    .O(\BAR0/BR-15-8/EQ3 )
  );
  X_INV   \NlwInverterBlock_BAR0/BR-15-8/X2/O  (
    .I(\NlwInverterSignal_BAR0/BR-15-8/X2/O ),
    .O(\BAR0/BR-15-8/EQ2 )
  );
  X_INV   \NlwInverterBlock_BAR0/BR-15-8/X0/O  (
    .I(\NlwInverterSignal_BAR0/BR-15-8/X0/O ),
    .O(\BAR0/BR-15-8/EQ0 )
  );
  X_INV   \NlwInverterBlock_BAR0/BR-15-8/X4/O  (
    .I(\NlwInverterSignal_BAR0/BR-15-8/X4/O ),
    .O(\BAR0/BR-15-8/EQ4 )
  );
  X_INV   \NlwInverterBlock_BAR0/BR-15-8/X6/O  (
    .I(\NlwInverterSignal_BAR0/BR-15-8/X6/O ),
    .O(\BAR0/BR-15-8/EQ6 )
  );
  X_INV   \NlwInverterBlock_BAR0/BR-15-8/X7/O  (
    .I(\NlwInverterSignal_BAR0/BR-15-8/X7/O ),
    .O(\BAR0/BR-15-8/EQ7 )
  );
  X_INV   \NlwInverterBlock_BAR0/BR-15-8/X5/O  (
    .I(\NlwInverterSignal_BAR0/BR-15-8/X5/O ),
    .O(\BAR0/BR-15-8/EQ5 )
  );
  X_INV   \NlwInverterBlock_BAR0/BR-CMD/$1I194/I0  (
    .I(CBE_IN0),
    .O(\NlwInverterSignal_BAR0/BR-CMD/$1I194/I0 )
  );
  X_INV   \NlwInverterBlock_BAR0/BR-CMD/$1I173/I0  (
    .I(CBE_IN3),
    .O(\NlwInverterSignal_BAR0/BR-CMD/$1I173/I0 )
  );
  X_INV   \NlwInverterBlock_BAR0/BR-CMD/$1I173/I1  (
    .I(CBE_IN2),
    .O(\NlwInverterSignal_BAR0/BR-CMD/$1I173/I1 )
  );
  X_INV   \NlwInverterBlock_BAR0/BR-CMD/$1I117/I0  (
    .I(CFG36),
    .O(\NlwInverterSignal_BAR0/BR-CMD/$1I117/I0 )
  );
  X_INV   \NlwInverterBlock_BAR0/BR-CMD/$1I110/I0  (
    .I(CFG36),
    .O(\NlwInverterSignal_BAR0/BR-CMD/$1I110/I0 )
  );
  X_INV   \NlwInverterBlock_BAR0/BR-CMD/$1I100/I0  (
    .I(CFG36),
    .O(\NlwInverterSignal_BAR0/BR-CMD/$1I100/I0 )
  );
  X_INV   \NlwInverterBlock_BAR0/BR-CMD/$1I223/$1I31/I0  (
    .I(CFG36),
    .O(\NlwInverterSignal_BAR0/BR-CMD/$1I223/$1I31/I0 )
  );
  X_INV   \NlwInverterBlock_BAR0/BR-7-4/X7/O  (
    .I(\NlwInverterSignal_BAR0/BR-7-4/X7/O ),
    .O(\BAR0/BR-7-4/EQ7 )
  );
  X_INV   \NlwInverterBlock_BAR0/BR-7-4/X6/O  (
    .I(\NlwInverterSignal_BAR0/BR-7-4/X6/O ),
    .O(\BAR0/BR-7-4/EQ6 )
  );
  X_INV   \NlwInverterBlock_BAR0/BR-7-4/X5/O  (
    .I(\NlwInverterSignal_BAR0/BR-7-4/X5/O ),
    .O(\BAR0/BR-7-4/EQ5 )
  );
  X_INV   \NlwInverterBlock_BAR0/BR-7-4/X4/O  (
    .I(\NlwInverterSignal_BAR0/BR-7-4/X4/O ),
    .O(\BAR0/BR-7-4/EQ4 )
  );
  X_INV   \NlwInverterBlock_BAR0/$1I3440/$1I31/I0  (
    .I(CFG36),
    .O(\NlwInverterSignal_BAR0/$1I3440/$1I31/I0 )
  );
  X_INV   \NlwInverterBlock_BAR0/$1I3453/$1I31/I0  (
    .I(CFG36),
    .O(\NlwInverterSignal_BAR0/$1I3453/$1I31/I0 )
  );
  X_INV   \NlwInverterBlock_BAR0/$2I3321/$1I31/I0  (
    .I(CFG36),
    .O(\NlwInverterSignal_BAR0/$2I3321/$1I31/I0 )
  );
  X_INV   \NlwInverterBlock_BAR1/BR-31-24/X1/O  (
    .I(\NlwInverterSignal_BAR1/BR-31-24/X1/O ),
    .O(\BAR1/BR-31-24/EQ1 )
  );
  X_INV   \NlwInverterBlock_BAR1/BR-31-24/X3/O  (
    .I(\NlwInverterSignal_BAR1/BR-31-24/X3/O ),
    .O(\BAR1/BR-31-24/EQ3 )
  );
  X_INV   \NlwInverterBlock_BAR1/BR-31-24/X2/O  (
    .I(\NlwInverterSignal_BAR1/BR-31-24/X2/O ),
    .O(\BAR1/BR-31-24/EQ2 )
  );
  X_INV   \NlwInverterBlock_BAR1/BR-31-24/X0/O  (
    .I(\NlwInverterSignal_BAR1/BR-31-24/X0/O ),
    .O(\BAR1/BR-31-24/EQ0 )
  );
  X_INV   \NlwInverterBlock_BAR1/BR-31-24/X4/O  (
    .I(\NlwInverterSignal_BAR1/BR-31-24/X4/O ),
    .O(\BAR1/BR-31-24/EQ4 )
  );
  X_INV   \NlwInverterBlock_BAR1/BR-31-24/X6/O  (
    .I(\NlwInverterSignal_BAR1/BR-31-24/X6/O ),
    .O(\BAR1/BR-31-24/EQ6 )
  );
  X_INV   \NlwInverterBlock_BAR1/BR-31-24/X7/O  (
    .I(\NlwInverterSignal_BAR1/BR-31-24/X7/O ),
    .O(\BAR1/BR-31-24/EQ7 )
  );
  X_INV   \NlwInverterBlock_BAR1/BR-31-24/X5/O  (
    .I(\NlwInverterSignal_BAR1/BR-31-24/X5/O ),
    .O(\BAR1/BR-31-24/EQ5 )
  );
  X_INV   \NlwInverterBlock_BAR1/BR-23-16/X1/O  (
    .I(\NlwInverterSignal_BAR1/BR-23-16/X1/O ),
    .O(\BAR1/BR-23-16/EQ1 )
  );
  X_INV   \NlwInverterBlock_BAR1/BR-23-16/X3/O  (
    .I(\NlwInverterSignal_BAR1/BR-23-16/X3/O ),
    .O(\BAR1/BR-23-16/EQ3 )
  );
  X_INV   \NlwInverterBlock_BAR1/BR-23-16/X2/O  (
    .I(\NlwInverterSignal_BAR1/BR-23-16/X2/O ),
    .O(\BAR1/BR-23-16/EQ2 )
  );
  X_INV   \NlwInverterBlock_BAR1/BR-23-16/X0/O  (
    .I(\NlwInverterSignal_BAR1/BR-23-16/X0/O ),
    .O(\BAR1/BR-23-16/EQ0 )
  );
  X_INV   \NlwInverterBlock_BAR1/BR-23-16/X4/O  (
    .I(\NlwInverterSignal_BAR1/BR-23-16/X4/O ),
    .O(\BAR1/BR-23-16/EQ4 )
  );
  X_INV   \NlwInverterBlock_BAR1/BR-23-16/X6/O  (
    .I(\NlwInverterSignal_BAR1/BR-23-16/X6/O ),
    .O(\BAR1/BR-23-16/EQ6 )
  );
  X_INV   \NlwInverterBlock_BAR1/BR-23-16/X7/O  (
    .I(\NlwInverterSignal_BAR1/BR-23-16/X7/O ),
    .O(\BAR1/BR-23-16/EQ7 )
  );
  X_INV   \NlwInverterBlock_BAR1/BR-23-16/X5/O  (
    .I(\NlwInverterSignal_BAR1/BR-23-16/X5/O ),
    .O(\BAR1/BR-23-16/EQ5 )
  );
  X_INV   \NlwInverterBlock_BAR1/BR-15-8/X1/O  (
    .I(\NlwInverterSignal_BAR1/BR-15-8/X1/O ),
    .O(\BAR1/BR-15-8/EQ1 )
  );
  X_INV   \NlwInverterBlock_BAR1/BR-15-8/X3/O  (
    .I(\NlwInverterSignal_BAR1/BR-15-8/X3/O ),
    .O(\BAR1/BR-15-8/EQ3 )
  );
  X_INV   \NlwInverterBlock_BAR1/BR-15-8/X2/O  (
    .I(\NlwInverterSignal_BAR1/BR-15-8/X2/O ),
    .O(\BAR1/BR-15-8/EQ2 )
  );
  X_INV   \NlwInverterBlock_BAR1/BR-15-8/X0/O  (
    .I(\NlwInverterSignal_BAR1/BR-15-8/X0/O ),
    .O(\BAR1/BR-15-8/EQ0 )
  );
  X_INV   \NlwInverterBlock_BAR1/BR-15-8/X4/O  (
    .I(\NlwInverterSignal_BAR1/BR-15-8/X4/O ),
    .O(\BAR1/BR-15-8/EQ4 )
  );
  X_INV   \NlwInverterBlock_BAR1/BR-15-8/X6/O  (
    .I(\NlwInverterSignal_BAR1/BR-15-8/X6/O ),
    .O(\BAR1/BR-15-8/EQ6 )
  );
  X_INV   \NlwInverterBlock_BAR1/BR-15-8/X7/O  (
    .I(\NlwInverterSignal_BAR1/BR-15-8/X7/O ),
    .O(\BAR1/BR-15-8/EQ7 )
  );
  X_INV   \NlwInverterBlock_BAR1/BR-15-8/X5/O  (
    .I(\NlwInverterSignal_BAR1/BR-15-8/X5/O ),
    .O(\BAR1/BR-15-8/EQ5 )
  );
  X_INV   \NlwInverterBlock_BAR1/BR-CMD/$1I194/I0  (
    .I(CBE_IN0),
    .O(\NlwInverterSignal_BAR1/BR-CMD/$1I194/I0 )
  );
  X_INV   \NlwInverterBlock_BAR1/BR-CMD/$1I173/I0  (
    .I(CBE_IN3),
    .O(\NlwInverterSignal_BAR1/BR-CMD/$1I173/I0 )
  );
  X_INV   \NlwInverterBlock_BAR1/BR-CMD/$1I173/I1  (
    .I(CBE_IN2),
    .O(\NlwInverterSignal_BAR1/BR-CMD/$1I173/I1 )
  );
  X_INV   \NlwInverterBlock_BAR1/BR-CMD/$1I117/I0  (
    .I(CFG73),
    .O(\NlwInverterSignal_BAR1/BR-CMD/$1I117/I0 )
  );
  X_INV   \NlwInverterBlock_BAR1/BR-CMD/$1I110/I0  (
    .I(CFG73),
    .O(\NlwInverterSignal_BAR1/BR-CMD/$1I110/I0 )
  );
  X_INV   \NlwInverterBlock_BAR1/BR-CMD/$1I100/I0  (
    .I(CFG73),
    .O(\NlwInverterSignal_BAR1/BR-CMD/$1I100/I0 )
  );
  X_INV   \NlwInverterBlock_BAR1/BR-CMD/$1I223/$1I31/I0  (
    .I(CFG73),
    .O(\NlwInverterSignal_BAR1/BR-CMD/$1I223/$1I31/I0 )
  );
  X_INV   \NlwInverterBlock_BAR1/BR-7-4/X7/O  (
    .I(\NlwInverterSignal_BAR1/BR-7-4/X7/O ),
    .O(\BAR1/BR-7-4/EQ7 )
  );
  X_INV   \NlwInverterBlock_BAR1/BR-7-4/X6/O  (
    .I(\NlwInverterSignal_BAR1/BR-7-4/X6/O ),
    .O(\BAR1/BR-7-4/EQ6 )
  );
  X_INV   \NlwInverterBlock_BAR1/BR-7-4/X5/O  (
    .I(\NlwInverterSignal_BAR1/BR-7-4/X5/O ),
    .O(\BAR1/BR-7-4/EQ5 )
  );
  X_INV   \NlwInverterBlock_BAR1/BR-7-4/X4/O  (
    .I(\NlwInverterSignal_BAR1/BR-7-4/X4/O ),
    .O(\BAR1/BR-7-4/EQ4 )
  );
  X_INV   \NlwInverterBlock_BAR1/$1I3440/$1I31/I0  (
    .I(CFG73),
    .O(\NlwInverterSignal_BAR1/$1I3440/$1I31/I0 )
  );
  X_INV   \NlwInverterBlock_BAR1/$1I3453/$1I31/I0  (
    .I(CFG73),
    .O(\NlwInverterSignal_BAR1/$1I3453/$1I31/I0 )
  );
  X_INV   \NlwInverterBlock_BAR1/$2I3321/$1I31/I0  (
    .I(CFG73),
    .O(\NlwInverterSignal_BAR1/$2I3321/$1I31/I0 )
  );
  X_INV   \NlwInverterBlock_BAR2/BR-31-24/X1/O  (
    .I(\NlwInverterSignal_BAR2/BR-31-24/X1/O ),
    .O(\BAR2/BR-31-24/EQ1 )
  );
  X_INV   \NlwInverterBlock_BAR2/BR-31-24/X3/O  (
    .I(\NlwInverterSignal_BAR2/BR-31-24/X3/O ),
    .O(\BAR2/BR-31-24/EQ3 )
  );
  X_INV   \NlwInverterBlock_BAR2/BR-31-24/X2/O  (
    .I(\NlwInverterSignal_BAR2/BR-31-24/X2/O ),
    .O(\BAR2/BR-31-24/EQ2 )
  );
  X_INV   \NlwInverterBlock_BAR2/BR-31-24/X0/O  (
    .I(\NlwInverterSignal_BAR2/BR-31-24/X0/O ),
    .O(\BAR2/BR-31-24/EQ0 )
  );
  X_INV   \NlwInverterBlock_BAR2/BR-31-24/X4/O  (
    .I(\NlwInverterSignal_BAR2/BR-31-24/X4/O ),
    .O(\BAR2/BR-31-24/EQ4 )
  );
  X_INV   \NlwInverterBlock_BAR2/BR-31-24/X6/O  (
    .I(\NlwInverterSignal_BAR2/BR-31-24/X6/O ),
    .O(\BAR2/BR-31-24/EQ6 )
  );
  X_INV   \NlwInverterBlock_BAR2/BR-31-24/X7/O  (
    .I(\NlwInverterSignal_BAR2/BR-31-24/X7/O ),
    .O(\BAR2/BR-31-24/EQ7 )
  );
  X_INV   \NlwInverterBlock_BAR2/BR-31-24/X5/O  (
    .I(\NlwInverterSignal_BAR2/BR-31-24/X5/O ),
    .O(\BAR2/BR-31-24/EQ5 )
  );
  X_INV   \NlwInverterBlock_BAR2/BR-23-16/X1/O  (
    .I(\NlwInverterSignal_BAR2/BR-23-16/X1/O ),
    .O(\BAR2/BR-23-16/EQ1 )
  );
  X_INV   \NlwInverterBlock_BAR2/BR-23-16/X3/O  (
    .I(\NlwInverterSignal_BAR2/BR-23-16/X3/O ),
    .O(\BAR2/BR-23-16/EQ3 )
  );
  X_INV   \NlwInverterBlock_BAR2/BR-23-16/X2/O  (
    .I(\NlwInverterSignal_BAR2/BR-23-16/X2/O ),
    .O(\BAR2/BR-23-16/EQ2 )
  );
  X_INV   \NlwInverterBlock_BAR2/BR-23-16/X0/O  (
    .I(\NlwInverterSignal_BAR2/BR-23-16/X0/O ),
    .O(\BAR2/BR-23-16/EQ0 )
  );
  X_INV   \NlwInverterBlock_BAR2/BR-23-16/X4/O  (
    .I(\NlwInverterSignal_BAR2/BR-23-16/X4/O ),
    .O(\BAR2/BR-23-16/EQ4 )
  );
  X_INV   \NlwInverterBlock_BAR2/BR-23-16/X6/O  (
    .I(\NlwInverterSignal_BAR2/BR-23-16/X6/O ),
    .O(\BAR2/BR-23-16/EQ6 )
  );
  X_INV   \NlwInverterBlock_BAR2/BR-23-16/X7/O  (
    .I(\NlwInverterSignal_BAR2/BR-23-16/X7/O ),
    .O(\BAR2/BR-23-16/EQ7 )
  );
  X_INV   \NlwInverterBlock_BAR2/BR-23-16/X5/O  (
    .I(\NlwInverterSignal_BAR2/BR-23-16/X5/O ),
    .O(\BAR2/BR-23-16/EQ5 )
  );
  X_INV   \NlwInverterBlock_BAR2/BR-15-8/X1/O  (
    .I(\NlwInverterSignal_BAR2/BR-15-8/X1/O ),
    .O(\BAR2/BR-15-8/EQ1 )
  );
  X_INV   \NlwInverterBlock_BAR2/BR-15-8/X3/O  (
    .I(\NlwInverterSignal_BAR2/BR-15-8/X3/O ),
    .O(\BAR2/BR-15-8/EQ3 )
  );
  X_INV   \NlwInverterBlock_BAR2/BR-15-8/X2/O  (
    .I(\NlwInverterSignal_BAR2/BR-15-8/X2/O ),
    .O(\BAR2/BR-15-8/EQ2 )
  );
  X_INV   \NlwInverterBlock_BAR2/BR-15-8/X0/O  (
    .I(\NlwInverterSignal_BAR2/BR-15-8/X0/O ),
    .O(\BAR2/BR-15-8/EQ0 )
  );
  X_INV   \NlwInverterBlock_BAR2/BR-15-8/X4/O  (
    .I(\NlwInverterSignal_BAR2/BR-15-8/X4/O ),
    .O(\BAR2/BR-15-8/EQ4 )
  );
  X_INV   \NlwInverterBlock_BAR2/BR-15-8/X6/O  (
    .I(\NlwInverterSignal_BAR2/BR-15-8/X6/O ),
    .O(\BAR2/BR-15-8/EQ6 )
  );
  X_INV   \NlwInverterBlock_BAR2/BR-15-8/X7/O  (
    .I(\NlwInverterSignal_BAR2/BR-15-8/X7/O ),
    .O(\BAR2/BR-15-8/EQ7 )
  );
  X_INV   \NlwInverterBlock_BAR2/BR-15-8/X5/O  (
    .I(\NlwInverterSignal_BAR2/BR-15-8/X5/O ),
    .O(\BAR2/BR-15-8/EQ5 )
  );
  X_INV   \NlwInverterBlock_BAR2/BR-CMD/$1I194/I0  (
    .I(CBE_IN0),
    .O(\NlwInverterSignal_BAR2/BR-CMD/$1I194/I0 )
  );
  X_INV   \NlwInverterBlock_BAR2/BR-CMD/$1I173/I0  (
    .I(CBE_IN3),
    .O(\NlwInverterSignal_BAR2/BR-CMD/$1I173/I0 )
  );
  X_INV   \NlwInverterBlock_BAR2/BR-CMD/$1I173/I1  (
    .I(CBE_IN2),
    .O(\NlwInverterSignal_BAR2/BR-CMD/$1I173/I1 )
  );
  X_INV   \NlwInverterBlock_BAR2/BR-CMD/$1I117/I0  (
    .I(CFG110),
    .O(\NlwInverterSignal_BAR2/BR-CMD/$1I117/I0 )
  );
  X_INV   \NlwInverterBlock_BAR2/BR-CMD/$1I110/I0  (
    .I(CFG110),
    .O(\NlwInverterSignal_BAR2/BR-CMD/$1I110/I0 )
  );
  X_INV   \NlwInverterBlock_BAR2/BR-CMD/$1I100/I0  (
    .I(CFG110),
    .O(\NlwInverterSignal_BAR2/BR-CMD/$1I100/I0 )
  );
  X_INV   \NlwInverterBlock_BAR2/BR-CMD/$1I223/$1I31/I0  (
    .I(CFG110),
    .O(\NlwInverterSignal_BAR2/BR-CMD/$1I223/$1I31/I0 )
  );
  X_INV   \NlwInverterBlock_BAR2/BR-7-4/X7/O  (
    .I(\NlwInverterSignal_BAR2/BR-7-4/X7/O ),
    .O(\BAR2/BR-7-4/EQ7 )
  );
  X_INV   \NlwInverterBlock_BAR2/BR-7-4/X6/O  (
    .I(\NlwInverterSignal_BAR2/BR-7-4/X6/O ),
    .O(\BAR2/BR-7-4/EQ6 )
  );
  X_INV   \NlwInverterBlock_BAR2/BR-7-4/X5/O  (
    .I(\NlwInverterSignal_BAR2/BR-7-4/X5/O ),
    .O(\BAR2/BR-7-4/EQ5 )
  );
  X_INV   \NlwInverterBlock_BAR2/BR-7-4/X4/O  (
    .I(\NlwInverterSignal_BAR2/BR-7-4/X4/O ),
    .O(\BAR2/BR-7-4/EQ4 )
  );
  X_INV   \NlwInverterBlock_BAR2/$1I3440/$1I31/I0  (
    .I(CFG110),
    .O(\NlwInverterSignal_BAR2/$1I3440/$1I31/I0 )
  );
  X_INV   \NlwInverterBlock_BAR2/$1I3453/$1I31/I0  (
    .I(CFG110),
    .O(\NlwInverterSignal_BAR2/$1I3453/$1I31/I0 )
  );
  X_INV   \NlwInverterBlock_BAR2/$2I3321/$1I31/I0  (
    .I(CFG110),
    .O(\NlwInverterSignal_BAR2/$2I3321/$1I31/I0 )
  );
  X_INV   \NlwInverterBlock_F/UPPER/T0/T  (
    .I(OE15),
    .O(\NlwInverterSignal_F/UPPER/T0/T )
  );
  X_INV   \NlwInverterBlock_F/UPPER/T1/T  (
    .I(OE15),
    .O(\NlwInverterSignal_F/UPPER/T1/T )
  );
  X_INV   \NlwInverterBlock_F/UPPER/T2/T  (
    .I(OE15),
    .O(\NlwInverterSignal_F/UPPER/T2/T )
  );
  X_INV   \NlwInverterBlock_F/UPPER/T3/T  (
    .I(OE15),
    .O(\NlwInverterSignal_F/UPPER/T3/T )
  );
  X_INV   \NlwInverterBlock_F/UPPER/T4/T  (
    .I(OE15),
    .O(\NlwInverterSignal_F/UPPER/T4/T )
  );
  X_INV   \NlwInverterBlock_F/UPPER/T5/T  (
    .I(OE15),
    .O(\NlwInverterSignal_F/UPPER/T5/T )
  );
  X_INV   \NlwInverterBlock_F/UPPER/T6/T  (
    .I(OE15),
    .O(\NlwInverterSignal_F/UPPER/T6/T )
  );
  X_INV   \NlwInverterBlock_F/UPPER/T7/T  (
    .I(OE15),
    .O(\NlwInverterSignal_F/UPPER/T7/T )
  );
  X_INV   \NlwInverterBlock_F/UPPER/T8/T  (
    .I(OE15),
    .O(\NlwInverterSignal_F/UPPER/T8/T )
  );
  X_INV   \NlwInverterBlock_F/UPPER/T9/T  (
    .I(OE15),
    .O(\NlwInverterSignal_F/UPPER/T9/T )
  );
  X_INV   \NlwInverterBlock_F/UPPER/T10/T  (
    .I(OE15),
    .O(\NlwInverterSignal_F/UPPER/T10/T )
  );
  X_INV   \NlwInverterBlock_F/UPPER/T11/T  (
    .I(OE15),
    .O(\NlwInverterSignal_F/UPPER/T11/T )
  );
  X_INV   \NlwInverterBlock_F/UPPER/T12/T  (
    .I(OE15),
    .O(\NlwInverterSignal_F/UPPER/T12/T )
  );
  X_INV   \NlwInverterBlock_F/UPPER/T13/T  (
    .I(OE15),
    .O(\NlwInverterSignal_F/UPPER/T13/T )
  );
  X_INV   \NlwInverterBlock_F/UPPER/T14/T  (
    .I(OE15),
    .O(\NlwInverterSignal_F/UPPER/T14/T )
  );
  X_INV   \NlwInverterBlock_F/UPPER/T15/T  (
    .I(OE15),
    .O(\NlwInverterSignal_F/UPPER/T15/T )
  );
  X_INV   \NlwInverterBlock_F/LOWER/T0/T  (
    .I(OE15),
    .O(\NlwInverterSignal_F/LOWER/T0/T )
  );
  X_INV   \NlwInverterBlock_F/LOWER/T1/T  (
    .I(OE15),
    .O(\NlwInverterSignal_F/LOWER/T1/T )
  );
  X_INV   \NlwInverterBlock_F/LOWER/T2/T  (
    .I(OE15),
    .O(\NlwInverterSignal_F/LOWER/T2/T )
  );
  X_INV   \NlwInverterBlock_F/LOWER/T3/T  (
    .I(OE15),
    .O(\NlwInverterSignal_F/LOWER/T3/T )
  );
  X_INV   \NlwInverterBlock_F/LOWER/T4/T  (
    .I(OE15),
    .O(\NlwInverterSignal_F/LOWER/T4/T )
  );
  X_INV   \NlwInverterBlock_F/LOWER/T5/T  (
    .I(OE15),
    .O(\NlwInverterSignal_F/LOWER/T5/T )
  );
  X_INV   \NlwInverterBlock_F/LOWER/T6/T  (
    .I(OE15),
    .O(\NlwInverterSignal_F/LOWER/T6/T )
  );
  X_INV   \NlwInverterBlock_F/LOWER/T7/T  (
    .I(OE15),
    .O(\NlwInverterSignal_F/LOWER/T7/T )
  );
  X_INV   \NlwInverterBlock_F/LOWER/T8/T  (
    .I(OE15),
    .O(\NlwInverterSignal_F/LOWER/T8/T )
  );
  X_INV   \NlwInverterBlock_F/LOWER/T9/T  (
    .I(OE15),
    .O(\NlwInverterSignal_F/LOWER/T9/T )
  );
  X_INV   \NlwInverterBlock_F/LOWER/T10/T  (
    .I(OE15),
    .O(\NlwInverterSignal_F/LOWER/T10/T )
  );
  X_INV   \NlwInverterBlock_F/LOWER/T11/T  (
    .I(OE15),
    .O(\NlwInverterSignal_F/LOWER/T11/T )
  );
  X_INV   \NlwInverterBlock_F/LOWER/T12/T  (
    .I(OE15),
    .O(\NlwInverterSignal_F/LOWER/T12/T )
  );
  X_INV   \NlwInverterBlock_F/LOWER/T13/T  (
    .I(OE15),
    .O(\NlwInverterSignal_F/LOWER/T13/T )
  );
  X_INV   \NlwInverterBlock_F/LOWER/T14/T  (
    .I(OE15),
    .O(\NlwInverterSignal_F/LOWER/T14/T )
  );
  X_INV   \NlwInverterBlock_F/LOWER/T15/T  (
    .I(OE15),
    .O(\NlwInverterSignal_F/LOWER/T15/T )
  );
  X_INV   \NlwInverterBlock_1/UPPER/T0/T  (
    .I(OE1),
    .O(\NlwInverterSignal_1/UPPER/T0/T )
  );
  X_INV   \NlwInverterBlock_1/UPPER/T1/T  (
    .I(OE1),
    .O(\NlwInverterSignal_1/UPPER/T1/T )
  );
  X_INV   \NlwInverterBlock_1/UPPER/T2/T  (
    .I(OE1),
    .O(\NlwInverterSignal_1/UPPER/T2/T )
  );
  X_INV   \NlwInverterBlock_1/UPPER/T3/T  (
    .I(OE1),
    .O(\NlwInverterSignal_1/UPPER/T3/T )
  );
  X_INV   \NlwInverterBlock_1/UPPER/T4/T  (
    .I(OE1),
    .O(\NlwInverterSignal_1/UPPER/T4/T )
  );
  X_INV   \NlwInverterBlock_1/UPPER/T5/T  (
    .I(OE1),
    .O(\NlwInverterSignal_1/UPPER/T5/T )
  );
  X_INV   \NlwInverterBlock_1/UPPER/T6/T  (
    .I(OE1),
    .O(\NlwInverterSignal_1/UPPER/T6/T )
  );
  X_INV   \NlwInverterBlock_1/UPPER/T7/T  (
    .I(OE1),
    .O(\NlwInverterSignal_1/UPPER/T7/T )
  );
  X_INV   \NlwInverterBlock_1/UPPER/T8/T  (
    .I(OE1),
    .O(\NlwInverterSignal_1/UPPER/T8/T )
  );
  X_INV   \NlwInverterBlock_1/UPPER/T9/T  (
    .I(OE1),
    .O(\NlwInverterSignal_1/UPPER/T9/T )
  );
  X_INV   \NlwInverterBlock_1/UPPER/T10/T  (
    .I(OE1),
    .O(\NlwInverterSignal_1/UPPER/T10/T )
  );
  X_INV   \NlwInverterBlock_1/UPPER/T11/T  (
    .I(OE1),
    .O(\NlwInverterSignal_1/UPPER/T11/T )
  );
  X_INV   \NlwInverterBlock_1/UPPER/T12/T  (
    .I(OE1),
    .O(\NlwInverterSignal_1/UPPER/T12/T )
  );
  X_INV   \NlwInverterBlock_1/UPPER/T13/T  (
    .I(OE1),
    .O(\NlwInverterSignal_1/UPPER/T13/T )
  );
  X_INV   \NlwInverterBlock_1/UPPER/T14/T  (
    .I(OE1),
    .O(\NlwInverterSignal_1/UPPER/T14/T )
  );
  X_INV   \NlwInverterBlock_1/UPPER/T15/T  (
    .I(OE1),
    .O(\NlwInverterSignal_1/UPPER/T15/T )
  );
  X_INV   \NlwInverterBlock_1/LOWER/T0/T  (
    .I(OE1),
    .O(\NlwInverterSignal_1/LOWER/T0/T )
  );
  X_INV   \NlwInverterBlock_1/LOWER/T1/T  (
    .I(OE1),
    .O(\NlwInverterSignal_1/LOWER/T1/T )
  );
  X_INV   \NlwInverterBlock_1/LOWER/T2/T  (
    .I(OE1),
    .O(\NlwInverterSignal_1/LOWER/T2/T )
  );
  X_INV   \NlwInverterBlock_1/LOWER/T3/T  (
    .I(OE1),
    .O(\NlwInverterSignal_1/LOWER/T3/T )
  );
  X_INV   \NlwInverterBlock_1/LOWER/T4/T  (
    .I(OE1),
    .O(\NlwInverterSignal_1/LOWER/T4/T )
  );
  X_INV   \NlwInverterBlock_1/LOWER/T5/T  (
    .I(OE1),
    .O(\NlwInverterSignal_1/LOWER/T5/T )
  );
  X_INV   \NlwInverterBlock_1/LOWER/T6/T  (
    .I(OE1),
    .O(\NlwInverterSignal_1/LOWER/T6/T )
  );
  X_INV   \NlwInverterBlock_1/LOWER/T7/T  (
    .I(OE1),
    .O(\NlwInverterSignal_1/LOWER/T7/T )
  );
  X_INV   \NlwInverterBlock_1/LOWER/T8/T  (
    .I(OE1),
    .O(\NlwInverterSignal_1/LOWER/T8/T )
  );
  X_INV   \NlwInverterBlock_1/LOWER/T9/T  (
    .I(OE1),
    .O(\NlwInverterSignal_1/LOWER/T9/T )
  );
  X_INV   \NlwInverterBlock_1/LOWER/T10/T  (
    .I(OE1),
    .O(\NlwInverterSignal_1/LOWER/T10/T )
  );
  X_INV   \NlwInverterBlock_1/LOWER/T11/T  (
    .I(OE1),
    .O(\NlwInverterSignal_1/LOWER/T11/T )
  );
  X_INV   \NlwInverterBlock_1/LOWER/T12/T  (
    .I(OE1),
    .O(\NlwInverterSignal_1/LOWER/T12/T )
  );
  X_INV   \NlwInverterBlock_1/LOWER/T13/T  (
    .I(OE1),
    .O(\NlwInverterSignal_1/LOWER/T13/T )
  );
  X_INV   \NlwInverterBlock_1/LOWER/T14/T  (
    .I(OE1),
    .O(\NlwInverterSignal_1/LOWER/T14/T )
  );
  X_INV   \NlwInverterBlock_1/LOWER/T15/T  (
    .I(OE1),
    .O(\NlwInverterSignal_1/LOWER/T15/T )
  );
  X_INV   \NlwInverterBlock_0/UPPER/T0/T  (
    .I(OE_ROM),
    .O(\NlwInverterSignal_0/UPPER/T0/T )
  );
  X_INV   \NlwInverterBlock_0/UPPER/T1/T  (
    .I(OE_ROM),
    .O(\NlwInverterSignal_0/UPPER/T1/T )
  );
  X_INV   \NlwInverterBlock_0/UPPER/T2/T  (
    .I(OE_ROM),
    .O(\NlwInverterSignal_0/UPPER/T2/T )
  );
  X_INV   \NlwInverterBlock_0/UPPER/T3/T  (
    .I(OE_ROM),
    .O(\NlwInverterSignal_0/UPPER/T3/T )
  );
  X_INV   \NlwInverterBlock_0/UPPER/T4/T  (
    .I(OE_ROM),
    .O(\NlwInverterSignal_0/UPPER/T4/T )
  );
  X_INV   \NlwInverterBlock_0/UPPER/T5/T  (
    .I(OE_ROM),
    .O(\NlwInverterSignal_0/UPPER/T5/T )
  );
  X_INV   \NlwInverterBlock_0/UPPER/T6/T  (
    .I(OE_ROM),
    .O(\NlwInverterSignal_0/UPPER/T6/T )
  );
  X_INV   \NlwInverterBlock_0/UPPER/T7/T  (
    .I(OE_ROM),
    .O(\NlwInverterSignal_0/UPPER/T7/T )
  );
  X_INV   \NlwInverterBlock_0/UPPER/T8/T  (
    .I(OE_ROM),
    .O(\NlwInverterSignal_0/UPPER/T8/T )
  );
  X_INV   \NlwInverterBlock_0/UPPER/T9/T  (
    .I(OE_ROM),
    .O(\NlwInverterSignal_0/UPPER/T9/T )
  );
  X_INV   \NlwInverterBlock_0/UPPER/T10/T  (
    .I(OE_ROM),
    .O(\NlwInverterSignal_0/UPPER/T10/T )
  );
  X_INV   \NlwInverterBlock_0/UPPER/T11/T  (
    .I(OE_ROM),
    .O(\NlwInverterSignal_0/UPPER/T11/T )
  );
  X_INV   \NlwInverterBlock_0/UPPER/T12/T  (
    .I(OE_ROM),
    .O(\NlwInverterSignal_0/UPPER/T12/T )
  );
  X_INV   \NlwInverterBlock_0/UPPER/T13/T  (
    .I(OE_ROM),
    .O(\NlwInverterSignal_0/UPPER/T13/T )
  );
  X_INV   \NlwInverterBlock_0/UPPER/T14/T  (
    .I(OE_ROM),
    .O(\NlwInverterSignal_0/UPPER/T14/T )
  );
  X_INV   \NlwInverterBlock_0/UPPER/T15/T  (
    .I(OE_ROM),
    .O(\NlwInverterSignal_0/UPPER/T15/T )
  );
  X_INV   \NlwInverterBlock_0/LOWER/T0/T  (
    .I(OE_ROM),
    .O(\NlwInverterSignal_0/LOWER/T0/T )
  );
  X_INV   \NlwInverterBlock_0/LOWER/T1/T  (
    .I(OE_ROM),
    .O(\NlwInverterSignal_0/LOWER/T1/T )
  );
  X_INV   \NlwInverterBlock_0/LOWER/T2/T  (
    .I(OE_ROM),
    .O(\NlwInverterSignal_0/LOWER/T2/T )
  );
  X_INV   \NlwInverterBlock_0/LOWER/T3/T  (
    .I(OE_ROM),
    .O(\NlwInverterSignal_0/LOWER/T3/T )
  );
  X_INV   \NlwInverterBlock_0/LOWER/T4/T  (
    .I(OE_ROM),
    .O(\NlwInverterSignal_0/LOWER/T4/T )
  );
  X_INV   \NlwInverterBlock_0/LOWER/T5/T  (
    .I(OE_ROM),
    .O(\NlwInverterSignal_0/LOWER/T5/T )
  );
  X_INV   \NlwInverterBlock_0/LOWER/T6/T  (
    .I(OE_ROM),
    .O(\NlwInverterSignal_0/LOWER/T6/T )
  );
  X_INV   \NlwInverterBlock_0/LOWER/T7/T  (
    .I(OE_ROM),
    .O(\NlwInverterSignal_0/LOWER/T7/T )
  );
  X_INV   \NlwInverterBlock_0/LOWER/T8/T  (
    .I(OE_ROM),
    .O(\NlwInverterSignal_0/LOWER/T8/T )
  );
  X_INV   \NlwInverterBlock_0/LOWER/T9/T  (
    .I(OE_ROM),
    .O(\NlwInverterSignal_0/LOWER/T9/T )
  );
  X_INV   \NlwInverterBlock_0/LOWER/T10/T  (
    .I(OE_ROM),
    .O(\NlwInverterSignal_0/LOWER/T10/T )
  );
  X_INV   \NlwInverterBlock_0/LOWER/T11/T  (
    .I(OE_ROM),
    .O(\NlwInverterSignal_0/LOWER/T11/T )
  );
  X_INV   \NlwInverterBlock_0/LOWER/T12/T  (
    .I(OE_ROM),
    .O(\NlwInverterSignal_0/LOWER/T12/T )
  );
  X_INV   \NlwInverterBlock_0/LOWER/T13/T  (
    .I(OE_ROM),
    .O(\NlwInverterSignal_0/LOWER/T13/T )
  );
  X_INV   \NlwInverterBlock_0/LOWER/T14/T  (
    .I(OE_ROM),
    .O(\NlwInverterSignal_0/LOWER/T14/T )
  );
  X_INV   \NlwInverterBlock_0/LOWER/T15/T  (
    .I(OE_ROM),
    .O(\NlwInverterSignal_0/LOWER/T15/T )
  );
  X_INV   \NlwInverterBlock_PCI-CSR/STATREG/Q14/$1I2230/I0  (
    .I(ADIO30),
    .O(\NlwInverterSignal_PCI-CSR/STATREG/Q14/$1I2230/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CSR/STATREG/Q14/$1I2233/$1I7/I0  (
    .I(CE1_3),
    .O(\NlwInverterSignal_PCI-CSR/STATREG/Q14/$1I2233/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CSR/STATREG/Q12/$1I2230/I0  (
    .I(ADIO28),
    .O(\NlwInverterSignal_PCI-CSR/STATREG/Q12/$1I2230/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CSR/STATREG/Q12/$1I2233/$1I7/I0  (
    .I(CE1_3),
    .O(\NlwInverterSignal_PCI-CSR/STATREG/Q12/$1I2233/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CSR/STATREG/Q8/$1I2230/I0  (
    .I(ADIO24),
    .O(\NlwInverterSignal_PCI-CSR/STATREG/Q8/$1I2230/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CSR/STATREG/Q8/$1I2233/$1I7/I0  (
    .I(CE1_3),
    .O(\NlwInverterSignal_PCI-CSR/STATREG/Q8/$1I2233/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CSR/STATREG/Q11/$1I2230/I0  (
    .I(ADIO27),
    .O(\NlwInverterSignal_PCI-CSR/STATREG/Q11/$1I2230/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CSR/STATREG/Q11/$1I2233/$1I7/I0  (
    .I(CE1_3),
    .O(\NlwInverterSignal_PCI-CSR/STATREG/Q11/$1I2233/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CSR/STATREG/Q13/$1I2230/I0  (
    .I(ADIO29),
    .O(\NlwInverterSignal_PCI-CSR/STATREG/Q13/$1I2230/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CSR/STATREG/Q13/$1I2233/$1I7/I0  (
    .I(CE1_3),
    .O(\NlwInverterSignal_PCI-CSR/STATREG/Q13/$1I2233/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CSR/STATREG/Q15/$1I2230/I0  (
    .I(ADIO31),
    .O(\NlwInverterSignal_PCI-CSR/STATREG/Q15/$1I2230/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CSR/STATREG/Q15/$1I2233/$1I7/I0  (
    .I(CE1_3),
    .O(\NlwInverterSignal_PCI-CSR/STATREG/Q15/$1I2233/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-ROM/$1I8330/I0  (
    .I(NlwRenamedSig_OI_ADDR7),
    .O(\NlwInverterSignal_PCI-ROM/$1I8330/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-ROM/$1I8330/I1  (
    .I(NlwRenamedSig_OI_ADDR6),
    .O(\NlwInverterSignal_PCI-ROM/$1I8330/I1 )
  );
  X_INV   \NlwInverterBlock_PCI-ROM/$1I8282/I0  (
    .I(NlwRenamedSig_OI_ADDR7),
    .O(\NlwInverterSignal_PCI-ROM/$1I8282/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-ROM/$1I8282/I1  (
    .I(NlwRenamedSig_OI_ADDR6),
    .O(\NlwInverterSignal_PCI-ROM/$1I8282/I1 )
  );
  X_INV   \NlwInverterBlock_PCI-ROM/$1I8282/I2  (
    .I(CFG114),
    .O(\NlwInverterSignal_PCI-ROM/$1I8282/I2 )
  );
  X_INV   \NlwInverterBlock_PCI-ROM/$1I8237/I0  (
    .I(NlwRenamedSig_OI_ADDR7),
    .O(\NlwInverterSignal_PCI-ROM/$1I8237/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-ROM/$1I8237/I1  (
    .I(NlwRenamedSig_OI_ADDR6),
    .O(\NlwInverterSignal_PCI-ROM/$1I8237/I1 )
  );
  X_INV   \NlwInverterBlock_PCI-ROM/$1I8227/I0  (
    .I(NlwRenamedSig_OI_ADDR7),
    .O(\NlwInverterSignal_PCI-ROM/$1I8227/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-ROM/$1I8227/I1  (
    .I(NlwRenamedSig_OI_ADDR6),
    .O(\NlwInverterSignal_PCI-ROM/$1I8227/I1 )
  );
  X_INV   \NlwInverterBlock_PCI-ROM/$1I8227/I2  (
    .I(CFG114),
    .O(\NlwInverterSignal_PCI-ROM/$1I8227/I2 )
  );
  X_INV   \NlwInverterBlock_PCI-ROM/$1I8110/I0  (
    .I(NlwRenamedSig_OI_ADDR7),
    .O(\NlwInverterSignal_PCI-ROM/$1I8110/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-ROM/$1I8110/I1  (
    .I(NlwRenamedSig_OI_ADDR6),
    .O(\NlwInverterSignal_PCI-ROM/$1I8110/I1 )
  );
  X_INV   \NlwInverterBlock_PCI-ROM/$1I8078/I0  (
    .I(NlwRenamedSig_OI_ADDR7),
    .O(\NlwInverterSignal_PCI-ROM/$1I8078/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-ROM/$1I8078/I1  (
    .I(NlwRenamedSig_OI_ADDR6),
    .O(\NlwInverterSignal_PCI-ROM/$1I8078/I1 )
  );
  X_INV   \NlwInverterBlock_$4I4029/$1I2610/$1I43/$1I30/$1I7/I0  (
    .I(\$4I4029/$1I2610/$1N48 ),
    .O(\NlwInverterSignal_$4I4029/$1I2610/$1I43/$1I30/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$4I4029/$1I2610/$1I53/$1I30/$1I7/I0  (
    .I(\$4I4029/$1I2610/$1N51 ),
    .O(\NlwInverterSignal_$4I4029/$1I2610/$1I53/$1I30/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$4I4029/$1I2610/$1I58/$1I30/$1I7/I0  (
    .I(\$4I4029/$1I2610/$1N56 ),
    .O(\NlwInverterSignal_$4I4029/$1I2610/$1I58/$1I30/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$4I4029/$1I2610/$1I59/$1I30/$1I7/I0  (
    .I(\$4I4029/$1I2610/$1N61 ),
    .O(\NlwInverterSignal_$4I4029/$1I2610/$1I59/$1I30/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$4I4029/$1I2610/$1I68/$1I30/$1I7/I0  (
    .I(\$4I4029/$1I2610/$1N66 ),
    .O(\NlwInverterSignal_$4I4029/$1I2610/$1I68/$1I30/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$4I4029/$1I2610/$1I73/$1I30/$1I7/I0  (
    .I(\$4I4029/$1I2610/$1N71 ),
    .O(\NlwInverterSignal_$4I4029/$1I2610/$1I73/$1I30/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$4I4029/$1I2610/$1I79/$1I30/$1I7/I0  (
    .I(\$4I4029/$1I2610/$1N81 ),
    .O(\NlwInverterSignal_$4I4029/$1I2610/$1I79/$1I30/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$4I4029/$1I2610/$1I84/$1I30/$1I7/I0  (
    .I(\$4I4029/$1I2610/$1N86 ),
    .O(\NlwInverterSignal_$4I4029/$1I2610/$1I84/$1I30/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$4I4029/$1I2637/$1I43/$1I30/$1I7/I0  (
    .I(\$4I4029/$1I2637/$1N48 ),
    .O(\NlwInverterSignal_$4I4029/$1I2637/$1I43/$1I30/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$4I4029/$1I2637/$1I53/$1I30/$1I7/I0  (
    .I(\$4I4029/$1I2637/$1N51 ),
    .O(\NlwInverterSignal_$4I4029/$1I2637/$1I53/$1I30/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$4I4029/$1I2637/$1I58/$1I30/$1I7/I0  (
    .I(\$4I4029/$1I2637/$1N56 ),
    .O(\NlwInverterSignal_$4I4029/$1I2637/$1I58/$1I30/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$4I4029/$1I2637/$1I59/$1I30/$1I7/I0  (
    .I(\$4I4029/$1I2637/$1N61 ),
    .O(\NlwInverterSignal_$4I4029/$1I2637/$1I59/$1I30/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$4I4029/$1I2637/$1I68/$1I30/$1I7/I0  (
    .I(\$4I4029/$1I2637/$1N66 ),
    .O(\NlwInverterSignal_$4I4029/$1I2637/$1I68/$1I30/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$4I4029/$1I2637/$1I73/$1I30/$1I7/I0  (
    .I(\$4I4029/$1I2637/$1N71 ),
    .O(\NlwInverterSignal_$4I4029/$1I2637/$1I73/$1I30/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$4I4029/$1I2637/$1I79/$1I30/$1I7/I0  (
    .I(\$4I4029/$1I2637/$1N81 ),
    .O(\NlwInverterSignal_$4I4029/$1I2637/$1I79/$1I30/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$4I4029/$1I2637/$1I84/$1I30/$1I7/I0  (
    .I(\$4I4029/$1I2637/$1N86 ),
    .O(\NlwInverterSignal_$4I4029/$1I2637/$1I84/$1I30/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$4I4029/$1I2645/$1I43/$1I30/$1I7/I0  (
    .I(\$4I4029/$1I2645/$1N48 ),
    .O(\NlwInverterSignal_$4I4029/$1I2645/$1I43/$1I30/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$4I4029/$1I2645/$1I53/$1I30/$1I7/I0  (
    .I(\$4I4029/$1I2645/$1N51 ),
    .O(\NlwInverterSignal_$4I4029/$1I2645/$1I53/$1I30/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$4I4029/$1I2645/$1I58/$1I30/$1I7/I0  (
    .I(\$4I4029/$1I2645/$1N56 ),
    .O(\NlwInverterSignal_$4I4029/$1I2645/$1I58/$1I30/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$4I4029/$1I2645/$1I59/$1I30/$1I7/I0  (
    .I(\$4I4029/$1I2645/$1N61 ),
    .O(\NlwInverterSignal_$4I4029/$1I2645/$1I59/$1I30/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$4I4029/$1I2645/$1I68/$1I30/$1I7/I0  (
    .I(\$4I4029/$1I2645/$1N66 ),
    .O(\NlwInverterSignal_$4I4029/$1I2645/$1I68/$1I30/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$4I4029/$1I2645/$1I73/$1I30/$1I7/I0  (
    .I(\$4I4029/$1I2645/$1N71 ),
    .O(\NlwInverterSignal_$4I4029/$1I2645/$1I73/$1I30/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$4I4029/$1I2645/$1I79/$1I30/$1I7/I0  (
    .I(\$4I4029/$1I2645/$1N81 ),
    .O(\NlwInverterSignal_$4I4029/$1I2645/$1I79/$1I30/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$4I4029/$1I2645/$1I84/$1I30/$1I7/I0  (
    .I(\$4I4029/$1I2645/$1N86 ),
    .O(\NlwInverterSignal_$4I4029/$1I2645/$1I84/$1I30/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$4I4029/$1I2653/$1I43/$1I30/$1I7/I0  (
    .I(\$4I4029/$1I2653/$1N48 ),
    .O(\NlwInverterSignal_$4I4029/$1I2653/$1I43/$1I30/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$4I4029/$1I2653/$1I53/$1I30/$1I7/I0  (
    .I(\$4I4029/$1I2653/$1N51 ),
    .O(\NlwInverterSignal_$4I4029/$1I2653/$1I53/$1I30/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$4I4029/$1I2653/$1I58/$1I30/$1I7/I0  (
    .I(\$4I4029/$1I2653/$1N56 ),
    .O(\NlwInverterSignal_$4I4029/$1I2653/$1I58/$1I30/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$4I4029/$1I2653/$1I59/$1I30/$1I7/I0  (
    .I(\$4I4029/$1I2653/$1N61 ),
    .O(\NlwInverterSignal_$4I4029/$1I2653/$1I59/$1I30/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$4I4029/$1I2653/$1I68/$1I30/$1I7/I0  (
    .I(\$4I4029/$1I2653/$1N66 ),
    .O(\NlwInverterSignal_$4I4029/$1I2653/$1I68/$1I30/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$4I4029/$1I2653/$1I73/$1I30/$1I7/I0  (
    .I(\$4I4029/$1I2653/$1N71 ),
    .O(\NlwInverterSignal_$4I4029/$1I2653/$1I73/$1I30/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$4I4029/$1I2653/$1I79/$1I30/$1I7/I0  (
    .I(\$4I4029/$1I2653/$1N81 ),
    .O(\NlwInverterSignal_$4I4029/$1I2653/$1I79/$1I30/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$4I4029/$1I2653/$1I84/$1I30/$1I7/I0  (
    .I(\$4I4029/$1I2653/$1N86 ),
    .O(\NlwInverterSignal_$4I4029/$1I2653/$1I84/$1I30/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$4I4029/$1I2661/$1I43/$1I30/$1I7/I0  (
    .I(\$4I4029/$1I2661/$1N48 ),
    .O(\NlwInverterSignal_$4I4029/$1I2661/$1I43/$1I30/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$4I4029/$1I2661/$1I53/$1I30/$1I7/I0  (
    .I(\$4I4029/$1I2661/$1N51 ),
    .O(\NlwInverterSignal_$4I4029/$1I2661/$1I53/$1I30/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$4I4029/$1I2661/$1I58/$1I30/$1I7/I0  (
    .I(\$4I4029/$1I2661/$1N56 ),
    .O(\NlwInverterSignal_$4I4029/$1I2661/$1I58/$1I30/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$4I4029/$1I2661/$1I59/$1I30/$1I7/I0  (
    .I(\$4I4029/$1I2661/$1N61 ),
    .O(\NlwInverterSignal_$4I4029/$1I2661/$1I59/$1I30/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$4I4029/$1I2661/$1I68/$1I30/$1I7/I0  (
    .I(\$4I4029/$1I2661/$1N66 ),
    .O(\NlwInverterSignal_$4I4029/$1I2661/$1I68/$1I30/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$4I4029/$1I2661/$1I73/$1I30/$1I7/I0  (
    .I(\$4I4029/$1I2661/$1N71 ),
    .O(\NlwInverterSignal_$4I4029/$1I2661/$1I73/$1I30/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$4I4029/$1I2661/$1I79/$1I30/$1I7/I0  (
    .I(\$4I4029/$1I2661/$1N81 ),
    .O(\NlwInverterSignal_$4I4029/$1I2661/$1I79/$1I30/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$4I4029/$1I2661/$1I84/$1I30/$1I7/I0  (
    .I(\$4I4029/$1I2661/$1N86 ),
    .O(\NlwInverterSignal_$4I4029/$1I2661/$1I84/$1I30/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_E/UPPER/T0/T  (
    .I(OE_ADI),
    .O(\NlwInverterSignal_E/UPPER/T0/T )
  );
  X_INV   \NlwInverterBlock_E/UPPER/T1/T  (
    .I(OE_ADI),
    .O(\NlwInverterSignal_E/UPPER/T1/T )
  );
  X_INV   \NlwInverterBlock_E/UPPER/T2/T  (
    .I(OE_ADI),
    .O(\NlwInverterSignal_E/UPPER/T2/T )
  );
  X_INV   \NlwInverterBlock_E/UPPER/T3/T  (
    .I(OE_ADI),
    .O(\NlwInverterSignal_E/UPPER/T3/T )
  );
  X_INV   \NlwInverterBlock_E/UPPER/T4/T  (
    .I(OE_ADI),
    .O(\NlwInverterSignal_E/UPPER/T4/T )
  );
  X_INV   \NlwInverterBlock_E/UPPER/T5/T  (
    .I(OE_ADI),
    .O(\NlwInverterSignal_E/UPPER/T5/T )
  );
  X_INV   \NlwInverterBlock_E/UPPER/T6/T  (
    .I(OE_ADI),
    .O(\NlwInverterSignal_E/UPPER/T6/T )
  );
  X_INV   \NlwInverterBlock_E/UPPER/T7/T  (
    .I(OE_ADI),
    .O(\NlwInverterSignal_E/UPPER/T7/T )
  );
  X_INV   \NlwInverterBlock_E/UPPER/T8/T  (
    .I(OE_ADI),
    .O(\NlwInverterSignal_E/UPPER/T8/T )
  );
  X_INV   \NlwInverterBlock_E/UPPER/T9/T  (
    .I(OE_ADI),
    .O(\NlwInverterSignal_E/UPPER/T9/T )
  );
  X_INV   \NlwInverterBlock_E/UPPER/T10/T  (
    .I(OE_ADI),
    .O(\NlwInverterSignal_E/UPPER/T10/T )
  );
  X_INV   \NlwInverterBlock_E/UPPER/T11/T  (
    .I(OE_ADI),
    .O(\NlwInverterSignal_E/UPPER/T11/T )
  );
  X_INV   \NlwInverterBlock_E/UPPER/T12/T  (
    .I(OE_ADI),
    .O(\NlwInverterSignal_E/UPPER/T12/T )
  );
  X_INV   \NlwInverterBlock_E/UPPER/T13/T  (
    .I(OE_ADI),
    .O(\NlwInverterSignal_E/UPPER/T13/T )
  );
  X_INV   \NlwInverterBlock_E/UPPER/T14/T  (
    .I(OE_ADI),
    .O(\NlwInverterSignal_E/UPPER/T14/T )
  );
  X_INV   \NlwInverterBlock_E/UPPER/T15/T  (
    .I(OE_ADI),
    .O(\NlwInverterSignal_E/UPPER/T15/T )
  );
  X_INV   \NlwInverterBlock_E/LOWER/T0/T  (
    .I(OE_ADI),
    .O(\NlwInverterSignal_E/LOWER/T0/T )
  );
  X_INV   \NlwInverterBlock_E/LOWER/T1/T  (
    .I(OE_ADI),
    .O(\NlwInverterSignal_E/LOWER/T1/T )
  );
  X_INV   \NlwInverterBlock_E/LOWER/T2/T  (
    .I(OE_ADI),
    .O(\NlwInverterSignal_E/LOWER/T2/T )
  );
  X_INV   \NlwInverterBlock_E/LOWER/T3/T  (
    .I(OE_ADI),
    .O(\NlwInverterSignal_E/LOWER/T3/T )
  );
  X_INV   \NlwInverterBlock_E/LOWER/T4/T  (
    .I(OE_ADI),
    .O(\NlwInverterSignal_E/LOWER/T4/T )
  );
  X_INV   \NlwInverterBlock_E/LOWER/T5/T  (
    .I(OE_ADI),
    .O(\NlwInverterSignal_E/LOWER/T5/T )
  );
  X_INV   \NlwInverterBlock_E/LOWER/T6/T  (
    .I(OE_ADI),
    .O(\NlwInverterSignal_E/LOWER/T6/T )
  );
  X_INV   \NlwInverterBlock_E/LOWER/T7/T  (
    .I(OE_ADI),
    .O(\NlwInverterSignal_E/LOWER/T7/T )
  );
  X_INV   \NlwInverterBlock_E/LOWER/T8/T  (
    .I(OE_ADI),
    .O(\NlwInverterSignal_E/LOWER/T8/T )
  );
  X_INV   \NlwInverterBlock_E/LOWER/T9/T  (
    .I(OE_ADI),
    .O(\NlwInverterSignal_E/LOWER/T9/T )
  );
  X_INV   \NlwInverterBlock_E/LOWER/T10/T  (
    .I(OE_ADI),
    .O(\NlwInverterSignal_E/LOWER/T10/T )
  );
  X_INV   \NlwInverterBlock_E/LOWER/T11/T  (
    .I(OE_ADI),
    .O(\NlwInverterSignal_E/LOWER/T11/T )
  );
  X_INV   \NlwInverterBlock_E/LOWER/T12/T  (
    .I(OE_ADI),
    .O(\NlwInverterSignal_E/LOWER/T12/T )
  );
  X_INV   \NlwInverterBlock_E/LOWER/T13/T  (
    .I(OE_ADI),
    .O(\NlwInverterSignal_E/LOWER/T13/T )
  );
  X_INV   \NlwInverterBlock_E/LOWER/T14/T  (
    .I(OE_ADI),
    .O(\NlwInverterSignal_E/LOWER/T14/T )
  );
  X_INV   \NlwInverterBlock_E/LOWER/T15/T  (
    .I(OE_ADI),
    .O(\NlwInverterSignal_E/LOWER/T15/T )
  );
  X_INV   \NlwInverterBlock_E64/UPPER/T0/T  (
    .I(DP64_T),
    .O(\NlwInverterSignal_E64/UPPER/T0/T )
  );
  X_INV   \NlwInverterBlock_E64/UPPER/T1/T  (
    .I(DP64_T),
    .O(\NlwInverterSignal_E64/UPPER/T1/T )
  );
  X_INV   \NlwInverterBlock_E64/UPPER/T2/T  (
    .I(DP64_T),
    .O(\NlwInverterSignal_E64/UPPER/T2/T )
  );
  X_INV   \NlwInverterBlock_E64/UPPER/T3/T  (
    .I(DP64_T),
    .O(\NlwInverterSignal_E64/UPPER/T3/T )
  );
  X_INV   \NlwInverterBlock_E64/UPPER/T4/T  (
    .I(DP64_T),
    .O(\NlwInverterSignal_E64/UPPER/T4/T )
  );
  X_INV   \NlwInverterBlock_E64/UPPER/T5/T  (
    .I(DP64_T),
    .O(\NlwInverterSignal_E64/UPPER/T5/T )
  );
  X_INV   \NlwInverterBlock_E64/UPPER/T6/T  (
    .I(DP64_T),
    .O(\NlwInverterSignal_E64/UPPER/T6/T )
  );
  X_INV   \NlwInverterBlock_E64/UPPER/T7/T  (
    .I(DP64_T),
    .O(\NlwInverterSignal_E64/UPPER/T7/T )
  );
  X_INV   \NlwInverterBlock_E64/UPPER/T8/T  (
    .I(DP64_T),
    .O(\NlwInverterSignal_E64/UPPER/T8/T )
  );
  X_INV   \NlwInverterBlock_E64/UPPER/T9/T  (
    .I(DP64_T),
    .O(\NlwInverterSignal_E64/UPPER/T9/T )
  );
  X_INV   \NlwInverterBlock_E64/UPPER/T10/T  (
    .I(DP64_T),
    .O(\NlwInverterSignal_E64/UPPER/T10/T )
  );
  X_INV   \NlwInverterBlock_E64/UPPER/T11/T  (
    .I(DP64_T),
    .O(\NlwInverterSignal_E64/UPPER/T11/T )
  );
  X_INV   \NlwInverterBlock_E64/UPPER/T12/T  (
    .I(DP64_T),
    .O(\NlwInverterSignal_E64/UPPER/T12/T )
  );
  X_INV   \NlwInverterBlock_E64/UPPER/T13/T  (
    .I(DP64_T),
    .O(\NlwInverterSignal_E64/UPPER/T13/T )
  );
  X_INV   \NlwInverterBlock_E64/UPPER/T14/T  (
    .I(DP64_T),
    .O(\NlwInverterSignal_E64/UPPER/T14/T )
  );
  X_INV   \NlwInverterBlock_E64/UPPER/T15/T  (
    .I(DP64_T),
    .O(\NlwInverterSignal_E64/UPPER/T15/T )
  );
  X_INV   \NlwInverterBlock_E64/LOWER/T0/T  (
    .I(DP64_T),
    .O(\NlwInverterSignal_E64/LOWER/T0/T )
  );
  X_INV   \NlwInverterBlock_E64/LOWER/T1/T  (
    .I(DP64_T),
    .O(\NlwInverterSignal_E64/LOWER/T1/T )
  );
  X_INV   \NlwInverterBlock_E64/LOWER/T2/T  (
    .I(DP64_T),
    .O(\NlwInverterSignal_E64/LOWER/T2/T )
  );
  X_INV   \NlwInverterBlock_E64/LOWER/T3/T  (
    .I(DP64_T),
    .O(\NlwInverterSignal_E64/LOWER/T3/T )
  );
  X_INV   \NlwInverterBlock_E64/LOWER/T4/T  (
    .I(DP64_T),
    .O(\NlwInverterSignal_E64/LOWER/T4/T )
  );
  X_INV   \NlwInverterBlock_E64/LOWER/T5/T  (
    .I(DP64_T),
    .O(\NlwInverterSignal_E64/LOWER/T5/T )
  );
  X_INV   \NlwInverterBlock_E64/LOWER/T6/T  (
    .I(DP64_T),
    .O(\NlwInverterSignal_E64/LOWER/T6/T )
  );
  X_INV   \NlwInverterBlock_E64/LOWER/T7/T  (
    .I(DP64_T),
    .O(\NlwInverterSignal_E64/LOWER/T7/T )
  );
  X_INV   \NlwInverterBlock_E64/LOWER/T8/T  (
    .I(DP64_T),
    .O(\NlwInverterSignal_E64/LOWER/T8/T )
  );
  X_INV   \NlwInverterBlock_E64/LOWER/T9/T  (
    .I(DP64_T),
    .O(\NlwInverterSignal_E64/LOWER/T9/T )
  );
  X_INV   \NlwInverterBlock_E64/LOWER/T10/T  (
    .I(DP64_T),
    .O(\NlwInverterSignal_E64/LOWER/T10/T )
  );
  X_INV   \NlwInverterBlock_E64/LOWER/T11/T  (
    .I(DP64_T),
    .O(\NlwInverterSignal_E64/LOWER/T11/T )
  );
  X_INV   \NlwInverterBlock_E64/LOWER/T12/T  (
    .I(DP64_T),
    .O(\NlwInverterSignal_E64/LOWER/T12/T )
  );
  X_INV   \NlwInverterBlock_E64/LOWER/T13/T  (
    .I(DP64_T),
    .O(\NlwInverterSignal_E64/LOWER/T13/T )
  );
  X_INV   \NlwInverterBlock_E64/LOWER/T14/T  (
    .I(DP64_T),
    .O(\NlwInverterSignal_E64/LOWER/T14/T )
  );
  X_INV   \NlwInverterBlock_E64/LOWER/T15/T  (
    .I(DP64_T),
    .O(\NlwInverterSignal_E64/LOWER/T15/T )
  );
  X_INV   \NlwInverterBlock_OEADI/$1I4041/I0  (
    .I(IDLE_DUP),
    .O(\NlwInverterSignal_OEADI/$1I4041/I0 )
  );
  X_INV   \NlwInverterBlock_OEADI/$1I4040/I0  (
    .I(\FRAME- ),
    .O(\NlwInverterSignal_OEADI/$1I4040/I0 )
  );
  X_INV   \NlwInverterBlock_OEADI/$1I4031/I0  (
    .I(OLDKEEPOUT),
    .O(\NlwInverterSignal_OEADI/$1I4031/I0 )
  );
  X_INV   \NlwInverterBlock_OEADI/$1I4031/I1  (
    .I(\OEADI/CFG_SELFQ ),
    .O(\NlwInverterSignal_OEADI/$1I4031/I1 )
  );
  X_INV   \NlwInverterBlock_OEADI/$1I4031/I2  (
    .I(M_WRDN),
    .O(\NlwInverterSignal_OEADI/$1I4031/I2 )
  );
  X_INV   \NlwInverterBlock_OEADI/$1I4031/O  (
    .I(\NlwInverterSignal_OEADI/$1I4031/O ),
    .O(\OEADI/OAI64_0 )
  );
  X_INV   \NlwInverterBlock_OEADI/$1I4028/I0  (
    .I(\OEADI/MIDDLE ),
    .O(\NlwInverterSignal_OEADI/$1I4028/I0 )
  );
  X_INV   \NlwInverterBlock_OEADI/$1I4028/O  (
    .I(\NlwInverterSignal_OEADI/$1I4028/O ),
    .O(\OEADI/OAI64_1 )
  );
  X_INV   \NlwInverterBlock_OEADI/$1I3984/I0  (
    .I(\OEADI/MIDDLE ),
    .O(\NlwInverterSignal_OEADI/$1I3984/I0 )
  );
  X_INV   \NlwInverterBlock_OEADI/$1I3984/O  (
    .I(\NlwInverterSignal_OEADI/$1I3984/O ),
    .O(\OEADI/OAI32_1 )
  );
  X_INV   \NlwInverterBlock_OEADI/$1I3954/I0  (
    .I(OLDKEEPOUT),
    .O(\NlwInverterSignal_OEADI/$1I3954/I0 )
  );
  X_INV   \NlwInverterBlock_OEADI/$1I3954/I1  (
    .I(\OEADI/CFG_SELFQ ),
    .O(\NlwInverterSignal_OEADI/$1I3954/I1 )
  );
  X_INV   \NlwInverterBlock_OEADI/$1I3954/I2  (
    .I(M_WRDN),
    .O(\NlwInverterSignal_OEADI/$1I3954/I2 )
  );
  X_INV   \NlwInverterBlock_OEADI/$1I3954/O  (
    .I(\NlwInverterSignal_OEADI/$1I3954/O ),
    .O(\OEADI/OAI32_0 )
  );
  X_INV   \NlwInverterBlock_OEADI/$1I3864/I0  (
    .I(\FRAME- ),
    .O(\NlwInverterSignal_OEADI/$1I3864/I0 )
  );
  X_INV   \NlwInverterBlock_OEADI/$1I3860/I0  (
    .I(IDLE_DUP),
    .O(\NlwInverterSignal_OEADI/$1I3860/I0 )
  );
  X_INV   \NlwInverterBlock_$5I3771/$1I7/I0  (
    .I(CFG111),
    .O(\NlwInverterSignal_$5I3771/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$5I3781/$1I7/I0  (
    .I(CFG111),
    .O(\NlwInverterSignal_$5I3781/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_DEVSEL/$1I2310/M01/$1I31/I0  (
    .I(CFG247),
    .O(\NlwInverterSignal_DEVSEL/$1I2310/M01/$1I31/I0 )
  );
  X_INV   \NlwInverterBlock_DEVSEL/$1I2310/M23/$1I31/I0  (
    .I(CFG247),
    .O(\NlwInverterSignal_DEVSEL/$1I2310/M23/$1I31/I0 )
  );
  X_INV   \NlwInverterBlock_ACK64/$1I2310/M01/$1I31/I0  (
    .I(CFG247),
    .O(\NlwInverterSignal_ACK64/$1I2310/M01/$1I31/I0 )
  );
  X_INV   \NlwInverterBlock_ACK64/$1I2310/M23/$1I31/I0  (
    .I(CFG247),
    .O(\NlwInverterSignal_ACK64/$1I2310/M23/$1I31/I0 )
  );
  X_INV   \NlwInverterBlock_FRAME/$1I2310/M01/$1I31/I0  (
    .I(CFG247),
    .O(\NlwInverterSignal_FRAME/$1I2310/M01/$1I31/I0 )
  );
  X_INV   \NlwInverterBlock_FRAME/$1I2310/M23/$1I31/I0  (
    .I(CFG247),
    .O(\NlwInverterSignal_FRAME/$1I2310/M23/$1I31/I0 )
  );
  X_INV   \NlwInverterBlock_TRDY/$1I2310/M01/$1I31/I0  (
    .I(CFG247),
    .O(\NlwInverterSignal_TRDY/$1I2310/M01/$1I31/I0 )
  );
  X_INV   \NlwInverterBlock_TRDY/$1I2310/M23/$1I31/I0  (
    .I(CFG247),
    .O(\NlwInverterSignal_TRDY/$1I2310/M23/$1I31/I0 )
  );
  X_INV   \NlwInverterBlock_REQ64/$1I2310/M01/$1I31/I0  (
    .I(CFG247),
    .O(\NlwInverterSignal_REQ64/$1I2310/M01/$1I31/I0 )
  );
  X_INV   \NlwInverterBlock_REQ64/$1I2310/M23/$1I31/I0  (
    .I(CFG247),
    .O(\NlwInverterSignal_REQ64/$1I2310/M23/$1I31/I0 )
  );
  X_INV   \NlwInverterBlock_IRDY/$1I2310/M01/$1I31/I0  (
    .I(CFG247),
    .O(\NlwInverterSignal_IRDY/$1I2310/M01/$1I31/I0 )
  );
  X_INV   \NlwInverterBlock_IRDY/$1I2310/M23/$1I31/I0  (
    .I(CFG247),
    .O(\NlwInverterSignal_IRDY/$1I2310/M23/$1I31/I0 )
  );
  X_INV   \NlwInverterBlock_STOP/$1I2310/M01/$1I31/I0  (
    .I(CFG247),
    .O(\NlwInverterSignal_STOP/$1I2310/M01/$1I31/I0 )
  );
  X_INV   \NlwInverterBlock_STOP/$1I2310/M23/$1I31/I0  (
    .I(CFG247),
    .O(\NlwInverterSignal_STOP/$1I2310/M23/$1I31/I0 )
  );
  X_INV   \NlwInverterBlock_$7I576/$1I7/I0  (
    .I(CFG240),
    .O(\NlwInverterSignal_$7I576/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$7I577/$1I7/I0  (
    .I(CFG240),
    .O(\NlwInverterSignal_$7I577/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$7I622/$1I7/I0  (
    .I(CFG240),
    .O(\NlwInverterSignal_$7I622/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$7I623/$1I7/I0  (
    .I(CFG240),
    .O(\NlwInverterSignal_$7I623/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$7I824/$1I7/I0  (
    .I(CFG255),
    .O(\NlwInverterSignal_$7I824/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$7I826/$1I7/I0  (
    .I(CFG255),
    .O(\NlwInverterSignal_$7I826/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$7I828/$1I7/I0  (
    .I(CFG255),
    .O(\NlwInverterSignal_$7I828/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$7I830/$1I7/I0  (
    .I(CFG255),
    .O(\NlwInverterSignal_$7I830/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$7I832/$1I7/I0  (
    .I(CFG255),
    .O(\NlwInverterSignal_$7I832/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$7I834/$1I7/I0  (
    .I(CFG255),
    .O(\NlwInverterSignal_$7I834/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$7I836/$1I7/I0  (
    .I(CFG255),
    .O(\NlwInverterSignal_$7I836/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_$7I838/$1I7/I0  (
    .I(CFG255),
    .O(\NlwInverterSignal_$7I838/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CBE/$1I2773/I0  (
    .I(\IIRDY_I- ),
    .O(\NlwInverterSignal_PCI-CBE/$1I2773/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CBE/IO3/$1I2296/$1I7/I0  (
    .I(OUT_SEL),
    .O(\NlwInverterSignal_PCI-CBE/IO3/$1I2296/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CBE/IO3/$1I2303/$1I7/I0  (
    .I(\PCI-CBE/IO3/$1N2321 ),
    .O(\NlwInverterSignal_PCI-CBE/IO3/$1I2303/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CBE/IO2/$1I2296/$1I7/I0  (
    .I(OUT_SEL),
    .O(\NlwInverterSignal_PCI-CBE/IO2/$1I2296/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CBE/IO2/$1I2303/$1I7/I0  (
    .I(\PCI-CBE/IO2/$1N2321 ),
    .O(\NlwInverterSignal_PCI-CBE/IO2/$1I2303/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CBE/IO1/$1I2296/$1I7/I0  (
    .I(OUT_SEL),
    .O(\NlwInverterSignal_PCI-CBE/IO1/$1I2296/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CBE/IO1/$1I2303/$1I7/I0  (
    .I(\PCI-CBE/IO1/$1N2321 ),
    .O(\NlwInverterSignal_PCI-CBE/IO1/$1I2303/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CBE/IO0/$1I2296/$1I7/I0  (
    .I(OUT_SEL),
    .O(\NlwInverterSignal_PCI-CBE/IO0/$1I2296/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CBE/IO0/$1I2303/$1I7/I0  (
    .I(\PCI-CBE/IO0/$1N2321 ),
    .O(\NlwInverterSignal_PCI-CBE/IO0/$1I2303/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CBE/$1I2777/$1I7/I0  (
    .I(CFG253),
    .O(\NlwInverterSignal_PCI-CBE/$1I2777/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CBE/$1I2779/$1I7/I0  (
    .I(CFG253),
    .O(\NlwInverterSignal_PCI-CBE/$1I2779/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/IO28/$1I2246/$1I7/I0  (
    .I(FAIL64_INT),
    .O(\NlwInverterSignal_PCI-AD/IO28/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/IO30/$1I2246/$1I7/I0  (
    .I(FAIL64_INT),
    .O(\NlwInverterSignal_PCI-AD/IO30/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/IO29/$1I2246/$1I7/I0  (
    .I(FAIL64_INT),
    .O(\NlwInverterSignal_PCI-AD/IO29/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/IO31/$1I2246/$1I7/I0  (
    .I(FAIL64_INT),
    .O(\NlwInverterSignal_PCI-AD/IO31/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/IO20/$1I2246/$1I7/I0  (
    .I(FAIL64_INT),
    .O(\NlwInverterSignal_PCI-AD/IO20/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/IO22/$1I2246/$1I7/I0  (
    .I(FAIL64_INT),
    .O(\NlwInverterSignal_PCI-AD/IO22/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/IO21/$1I2246/$1I7/I0  (
    .I(FAIL64_INT),
    .O(\NlwInverterSignal_PCI-AD/IO21/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/IO23/$1I2246/$1I7/I0  (
    .I(FAIL64_INT),
    .O(\NlwInverterSignal_PCI-AD/IO23/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/IO12/$1I2246/$1I7/I0  (
    .I(FAIL64_INT),
    .O(\NlwInverterSignal_PCI-AD/IO12/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/IO14/$1I2246/$1I7/I0  (
    .I(FAIL64_INT),
    .O(\NlwInverterSignal_PCI-AD/IO14/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/IO13/$1I2246/$1I7/I0  (
    .I(FAIL64_INT),
    .O(\NlwInverterSignal_PCI-AD/IO13/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/IO15/$1I2246/$1I7/I0  (
    .I(FAIL64_INT),
    .O(\NlwInverterSignal_PCI-AD/IO15/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/IO4/$1I2246/$1I7/I0  (
    .I(FAIL64_INT),
    .O(\NlwInverterSignal_PCI-AD/IO4/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/IO6/$1I2246/$1I7/I0  (
    .I(FAIL64_INT),
    .O(\NlwInverterSignal_PCI-AD/IO6/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/IO5/$1I2246/$1I7/I0  (
    .I(FAIL64_INT),
    .O(\NlwInverterSignal_PCI-AD/IO5/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/IO7/$1I2246/$1I7/I0  (
    .I(FAIL64_INT),
    .O(\NlwInverterSignal_PCI-AD/IO7/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/$1I2927/$1I7/I0  (
    .I(OUT_SEL),
    .O(\NlwInverterSignal_PCI-AD/$1I2927/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/$1I2928/$1I7/I0  (
    .I(OUT_SEL),
    .O(\NlwInverterSignal_PCI-AD/$1I2928/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/$1I2929/$1I7/I0  (
    .I(OUT_SEL),
    .O(\NlwInverterSignal_PCI-AD/$1I2929/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/$1I2930/$1I7/I0  (
    .I(OUT_SEL),
    .O(\NlwInverterSignal_PCI-AD/$1I2930/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/$1I2931/$1I7/I0  (
    .I(OUT_SEL),
    .O(\NlwInverterSignal_PCI-AD/$1I2931/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/$1I2932/$1I7/I0  (
    .I(OUT_SEL),
    .O(\NlwInverterSignal_PCI-AD/$1I2932/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/$1I2933/$1I7/I0  (
    .I(OUT_SEL),
    .O(\NlwInverterSignal_PCI-AD/$1I2933/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/$1I2934/$1I7/I0  (
    .I(OUT_SEL),
    .O(\NlwInverterSignal_PCI-AD/$1I2934/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/$1I2935/$1I7/I0  (
    .I(OUT_SEL),
    .O(\NlwInverterSignal_PCI-AD/$1I2935/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/$1I2936/$1I7/I0  (
    .I(OUT_SEL),
    .O(\NlwInverterSignal_PCI-AD/$1I2936/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/$1I2937/$1I7/I0  (
    .I(OUT_SEL),
    .O(\NlwInverterSignal_PCI-AD/$1I2937/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/$1I2938/$1I7/I0  (
    .I(OUT_SEL),
    .O(\NlwInverterSignal_PCI-AD/$1I2938/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/$1I2939/$1I7/I0  (
    .I(OUT_SEL),
    .O(\NlwInverterSignal_PCI-AD/$1I2939/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/$1I2940/$1I7/I0  (
    .I(OUT_SEL),
    .O(\NlwInverterSignal_PCI-AD/$1I2940/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/$1I2941/$1I7/I0  (
    .I(OUT_SEL),
    .O(\NlwInverterSignal_PCI-AD/$1I2941/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/$1I2942/$1I7/I0  (
    .I(OUT_SEL),
    .O(\NlwInverterSignal_PCI-AD/$1I2942/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/$1I2943/$1I7/I0  (
    .I(OUT_SEL),
    .O(\NlwInverterSignal_PCI-AD/$1I2943/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/$1I2944/$1I7/I0  (
    .I(OUT_SEL),
    .O(\NlwInverterSignal_PCI-AD/$1I2944/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/$1I2945/$1I7/I0  (
    .I(OUT_SEL),
    .O(\NlwInverterSignal_PCI-AD/$1I2945/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/$1I2946/$1I7/I0  (
    .I(OUT_SEL),
    .O(\NlwInverterSignal_PCI-AD/$1I2946/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/$1I2947/$1I7/I0  (
    .I(OUT_SEL),
    .O(\NlwInverterSignal_PCI-AD/$1I2947/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/$1I2948/$1I7/I0  (
    .I(OUT_SEL),
    .O(\NlwInverterSignal_PCI-AD/$1I2948/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/$1I2949/$1I7/I0  (
    .I(OUT_SEL),
    .O(\NlwInverterSignal_PCI-AD/$1I2949/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/$1I2950/$1I7/I0  (
    .I(OUT_SEL),
    .O(\NlwInverterSignal_PCI-AD/$1I2950/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/$1I2951/$1I7/I0  (
    .I(OUT_SEL),
    .O(\NlwInverterSignal_PCI-AD/$1I2951/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/$1I2952/$1I7/I0  (
    .I(OUT_SEL),
    .O(\NlwInverterSignal_PCI-AD/$1I2952/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/$1I2953/$1I7/I0  (
    .I(OUT_SEL),
    .O(\NlwInverterSignal_PCI-AD/$1I2953/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/$1I2954/$1I7/I0  (
    .I(OUT_SEL),
    .O(\NlwInverterSignal_PCI-AD/$1I2954/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/$1I2955/$1I7/I0  (
    .I(OUT_SEL),
    .O(\NlwInverterSignal_PCI-AD/$1I2955/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/$1I2956/$1I7/I0  (
    .I(OUT_SEL),
    .O(\NlwInverterSignal_PCI-AD/$1I2956/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/$1I2957/$1I7/I0  (
    .I(OUT_SEL),
    .O(\NlwInverterSignal_PCI-AD/$1I2957/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/$1I2958/$1I7/I0  (
    .I(OUT_SEL),
    .O(\NlwInverterSignal_PCI-AD/$1I2958/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/IO27/$1I2246/$1I7/I0  (
    .I(FAIL64_INT),
    .O(\NlwInverterSignal_PCI-AD/IO27/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/IO26/$1I2246/$1I7/I0  (
    .I(FAIL64_INT),
    .O(\NlwInverterSignal_PCI-AD/IO26/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/IO25/$1I2246/$1I7/I0  (
    .I(FAIL64_INT),
    .O(\NlwInverterSignal_PCI-AD/IO25/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/IO24/$1I2246/$1I7/I0  (
    .I(FAIL64_INT),
    .O(\NlwInverterSignal_PCI-AD/IO24/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/IO19/$1I2246/$1I7/I0  (
    .I(FAIL64_INT),
    .O(\NlwInverterSignal_PCI-AD/IO19/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/IO18/$1I2246/$1I7/I0  (
    .I(FAIL64_INT),
    .O(\NlwInverterSignal_PCI-AD/IO18/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/IO17/$1I2246/$1I7/I0  (
    .I(FAIL64_INT),
    .O(\NlwInverterSignal_PCI-AD/IO17/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/IO16/$1I2246/$1I7/I0  (
    .I(FAIL64_INT),
    .O(\NlwInverterSignal_PCI-AD/IO16/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/IO11/$1I2246/$1I7/I0  (
    .I(FAIL64_INT),
    .O(\NlwInverterSignal_PCI-AD/IO11/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/IO10/$1I2246/$1I7/I0  (
    .I(FAIL64_INT),
    .O(\NlwInverterSignal_PCI-AD/IO10/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/IO9/$1I2246/$1I7/I0  (
    .I(FAIL64_INT),
    .O(\NlwInverterSignal_PCI-AD/IO9/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/IO8/$1I2246/$1I7/I0  (
    .I(FAIL64_INT),
    .O(\NlwInverterSignal_PCI-AD/IO8/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/IO3/$1I2246/$1I7/I0  (
    .I(FAIL64_INT),
    .O(\NlwInverterSignal_PCI-AD/IO3/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/IO2/$1I2246/$1I7/I0  (
    .I(FAIL64_INT),
    .O(\NlwInverterSignal_PCI-AD/IO2/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/IO1/$1I2246/$1I7/I0  (
    .I(FAIL64_INT),
    .O(\NlwInverterSignal_PCI-AD/IO1/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD/IO0/$1I2246/$1I7/I0  (
    .I(FAIL64_INT),
    .O(\NlwInverterSignal_PCI-AD/IO0/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD64/IO28/$1I2246/$1I7/I0  (
    .I(OUT_SEL64),
    .O(\NlwInverterSignal_PCI-AD64/IO28/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD64/IO30/$1I2246/$1I7/I0  (
    .I(OUT_SEL64),
    .O(\NlwInverterSignal_PCI-AD64/IO30/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD64/IO29/$1I2246/$1I7/I0  (
    .I(OUT_SEL64),
    .O(\NlwInverterSignal_PCI-AD64/IO29/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD64/IO31/$1I2246/$1I7/I0  (
    .I(OUT_SEL64),
    .O(\NlwInverterSignal_PCI-AD64/IO31/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD64/IO20/$1I2246/$1I7/I0  (
    .I(OUT_SEL64),
    .O(\NlwInverterSignal_PCI-AD64/IO20/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD64/IO22/$1I2246/$1I7/I0  (
    .I(OUT_SEL64),
    .O(\NlwInverterSignal_PCI-AD64/IO22/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD64/IO21/$1I2246/$1I7/I0  (
    .I(OUT_SEL64),
    .O(\NlwInverterSignal_PCI-AD64/IO21/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD64/IO23/$1I2246/$1I7/I0  (
    .I(OUT_SEL64),
    .O(\NlwInverterSignal_PCI-AD64/IO23/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD64/IO12/$1I2246/$1I7/I0  (
    .I(OUT_SEL64),
    .O(\NlwInverterSignal_PCI-AD64/IO12/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD64/IO14/$1I2246/$1I7/I0  (
    .I(OUT_SEL64),
    .O(\NlwInverterSignal_PCI-AD64/IO14/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD64/IO13/$1I2246/$1I7/I0  (
    .I(OUT_SEL64),
    .O(\NlwInverterSignal_PCI-AD64/IO13/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD64/IO15/$1I2246/$1I7/I0  (
    .I(OUT_SEL64),
    .O(\NlwInverterSignal_PCI-AD64/IO15/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD64/IO4/$1I2246/$1I7/I0  (
    .I(OUT_SEL64),
    .O(\NlwInverterSignal_PCI-AD64/IO4/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD64/IO6/$1I2246/$1I7/I0  (
    .I(OUT_SEL64),
    .O(\NlwInverterSignal_PCI-AD64/IO6/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD64/IO5/$1I2246/$1I7/I0  (
    .I(OUT_SEL64),
    .O(\NlwInverterSignal_PCI-AD64/IO5/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD64/IO7/$1I2246/$1I7/I0  (
    .I(OUT_SEL64),
    .O(\NlwInverterSignal_PCI-AD64/IO7/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD64/IO27/$1I2246/$1I7/I0  (
    .I(OUT_SEL64),
    .O(\NlwInverterSignal_PCI-AD64/IO27/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD64/IO26/$1I2246/$1I7/I0  (
    .I(OUT_SEL64),
    .O(\NlwInverterSignal_PCI-AD64/IO26/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD64/IO25/$1I2246/$1I7/I0  (
    .I(OUT_SEL64),
    .O(\NlwInverterSignal_PCI-AD64/IO25/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD64/IO24/$1I2246/$1I7/I0  (
    .I(OUT_SEL64),
    .O(\NlwInverterSignal_PCI-AD64/IO24/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD64/IO19/$1I2246/$1I7/I0  (
    .I(OUT_SEL64),
    .O(\NlwInverterSignal_PCI-AD64/IO19/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD64/IO18/$1I2246/$1I7/I0  (
    .I(OUT_SEL64),
    .O(\NlwInverterSignal_PCI-AD64/IO18/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD64/IO17/$1I2246/$1I7/I0  (
    .I(OUT_SEL64),
    .O(\NlwInverterSignal_PCI-AD64/IO17/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD64/IO16/$1I2246/$1I7/I0  (
    .I(OUT_SEL64),
    .O(\NlwInverterSignal_PCI-AD64/IO16/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD64/IO11/$1I2246/$1I7/I0  (
    .I(OUT_SEL64),
    .O(\NlwInverterSignal_PCI-AD64/IO11/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD64/IO10/$1I2246/$1I7/I0  (
    .I(OUT_SEL64),
    .O(\NlwInverterSignal_PCI-AD64/IO10/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD64/IO9/$1I2246/$1I7/I0  (
    .I(OUT_SEL64),
    .O(\NlwInverterSignal_PCI-AD64/IO9/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD64/IO8/$1I2246/$1I7/I0  (
    .I(OUT_SEL64),
    .O(\NlwInverterSignal_PCI-AD64/IO8/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD64/IO3/$1I2246/$1I7/I0  (
    .I(OUT_SEL64),
    .O(\NlwInverterSignal_PCI-AD64/IO3/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD64/IO2/$1I2246/$1I7/I0  (
    .I(OUT_SEL64),
    .O(\NlwInverterSignal_PCI-AD64/IO2/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD64/IO1/$1I2246/$1I7/I0  (
    .I(OUT_SEL64),
    .O(\NlwInverterSignal_PCI-AD64/IO1/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-AD64/IO0/$1I2246/$1I7/I0  (
    .I(OUT_SEL64),
    .O(\NlwInverterSignal_PCI-AD64/IO0/$1I2246/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CBE64/IO3/$1I2296/$1I7/I0  (
    .I(OUT_SEL64),
    .O(\NlwInverterSignal_PCI-CBE64/IO3/$1I2296/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CBE64/IO3/$1I2303/$1I7/I0  (
    .I(\PCI-CBE64/IO3/$1N2321 ),
    .O(\NlwInverterSignal_PCI-CBE64/IO3/$1I2303/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CBE64/IO2/$1I2296/$1I7/I0  (
    .I(OUT_SEL64),
    .O(\NlwInverterSignal_PCI-CBE64/IO2/$1I2296/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CBE64/IO2/$1I2303/$1I7/I0  (
    .I(\PCI-CBE64/IO2/$1N2321 ),
    .O(\NlwInverterSignal_PCI-CBE64/IO2/$1I2303/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CBE64/IO1/$1I2296/$1I7/I0  (
    .I(OUT_SEL64),
    .O(\NlwInverterSignal_PCI-CBE64/IO1/$1I2296/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CBE64/IO1/$1I2303/$1I7/I0  (
    .I(\PCI-CBE64/IO1/$1N2321 ),
    .O(\NlwInverterSignal_PCI-CBE64/IO1/$1I2303/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CBE64/IO0/$1I2296/$1I7/I0  (
    .I(OUT_SEL64),
    .O(\NlwInverterSignal_PCI-CBE64/IO0/$1I2296/$1I7/I0 )
  );
  X_INV   \NlwInverterBlock_PCI-CBE64/IO0/$1I2303/$1I7/I0  (
    .I(\PCI-CBE64/IO0/$1N2321 ),
    .O(\NlwInverterSignal_PCI-CBE64/IO0/$1I2303/$1I7/I0 )
  );
// synthesis translate_on
endmodule
